//ytydla_vinp.sv

//---------------------------------------
// YTYDLA Vector Inner Product
//---------------------------------------

module ytydla_vinp(ytydla_core_clk,
                   ytydla_core_rst_n,
                   mem2vinp_a_0,
                   mem2vinp_a_1,
                   mem2vinp_a_2,
                   mem2vinp_a_3,
                   mem2vinp_a_4,
                   mem2vinp_a_5,
                   mem2vinp_a_6,
                   mem2vinp_a_7,
                   mem2vinp_a_8,
                   mem2vinp_a_9,
                   mem2vinp_a_10,
                   mem2vinp_a_11,
                   mem2vinp_a_12,
                   mem2vinp_a_13,
                   mem2vinp_a_14,
                   mem2vinp_a_15,
                   mem2vinp_a_16,
                   mem2vinp_a_17,
                   mem2vinp_a_18,
                   mem2vinp_a_19,
                   mem2vinp_a_20,
                   mem2vinp_a_21,
                   mem2vinp_a_22,
                   mem2vinp_a_23,
                   mem2vinp_a_24,
                   mem2vinp_a_25,
                   mem2vinp_a_26,
                   mem2vinp_a_27,
                   mem2vinp_a_28,
                   mem2vinp_a_29,
                   mem2vinp_a_30,
                   mem2vinp_a_31,
                   mem2vinp_a_32,
                   mem2vinp_a_33,
                   mem2vinp_a_34,
                   mem2vinp_a_35,
                   mem2vinp_a_36,
                   mem2vinp_a_37,
                   mem2vinp_a_38,
                   mem2vinp_a_39,
                   mem2vinp_a_40,
                   mem2vinp_a_41,
                   mem2vinp_a_42,
                   mem2vinp_a_43,
                   mem2vinp_a_44,
                   mem2vinp_a_45,
                   mem2vinp_a_46,
                   mem2vinp_a_47,
                   mem2vinp_a_48,
                   mem2vinp_a_49,
                   mem2vinp_a_50,
                   mem2vinp_a_51,
                   mem2vinp_a_52,
                   mem2vinp_a_53,
                   mem2vinp_a_54,
                   mem2vinp_a_55,
                   mem2vinp_a_56,
                   mem2vinp_a_57,
                   mem2vinp_a_58,
                   mem2vinp_a_59,
                   mem2vinp_a_60,
                   mem2vinp_a_61,
                   mem2vinp_a_62,
                   mem2vinp_a_63,
                   mem2vinp_b_0,
                   mem2vinp_b_1,
                   mem2vinp_b_2,
                   mem2vinp_b_3,
                   mem2vinp_b_4,
                   mem2vinp_b_5,
                   mem2vinp_b_6,
                   mem2vinp_b_7,
                   mem2vinp_b_8,
                   mem2vinp_b_9,
                   mem2vinp_b_10,
                   mem2vinp_b_11,
                   mem2vinp_b_12,
                   mem2vinp_b_13,
                   mem2vinp_b_14,
                   mem2vinp_b_15,
                   mem2vinp_b_16,
                   mem2vinp_b_17,
                   mem2vinp_b_18,
                   mem2vinp_b_19,
                   mem2vinp_b_20,
                   mem2vinp_b_21,
                   mem2vinp_b_22,
                   mem2vinp_b_23,
                   mem2vinp_b_24,
                   mem2vinp_b_25,
                   mem2vinp_b_26,
                   mem2vinp_b_27,
                   mem2vinp_b_28,
                   mem2vinp_b_29,
                   mem2vinp_b_30,
                   mem2vinp_b_31,
                   mem2vinp_b_32,
                   mem2vinp_b_33,
                   mem2vinp_b_34,
                   mem2vinp_b_35,
                   mem2vinp_b_36,
                   mem2vinp_b_37,
                   mem2vinp_b_38,
                   mem2vinp_b_39,
                   mem2vinp_b_40,
                   mem2vinp_b_41,
                   mem2vinp_b_42,
                   mem2vinp_b_43,
                   mem2vinp_b_44,
                   mem2vinp_b_45,
                   mem2vinp_b_46,
                   mem2vinp_b_47,
                   mem2vinp_b_48,
                   mem2vinp_b_49,
                   mem2vinp_b_50,
                   mem2vinp_b_51,
                   mem2vinp_b_52,
                   mem2vinp_b_53,
                   mem2vinp_b_54,
                   mem2vinp_b_55,
                   mem2vinp_b_56,
                   mem2vinp_b_57,
                   mem2vinp_b_58,
                   mem2vinp_b_59,
                   mem2vinp_b_60,
                   mem2vinp_b_61,
                   mem2vinp_b_62,
                   mem2vinp_b_63,
                   mem2vinp_size,
                   vinp2mem_result_0,
                   vinp2mem_result_1,
                   vinp2mem_result_2,
                   vinp2mem_result_3,
                   vinp2mem_result_4,
                   vinp2mem_result_5,
                   vinp2mem_result_6,
                   vinp2mem_result_7,
                   vinp2mem_result_8,
                   vinp2mem_result_9,
                   vinp2mem_result_10,
                   vinp2mem_result_11,
                   vinp2mem_result_12,
                   vinp2mem_result_13,
                   vinp2mem_result_14,
                   vinp2mem_result_15,
                   vinp2mem_result_16,
                   vinp2mem_result_17,
                   vinp2mem_result_18,
                   vinp2mem_result_19,
                   vinp2mem_result_20,
                   vinp2mem_result_21,
                   vinp2mem_result_22,
                   vinp2mem_result_23,
                   vinp2mem_result_24,
                   vinp2mem_result_25,
                   vinp2mem_result_26,
                   vinp2mem_result_27,
                   vinp2mem_result_28,
                   vinp2mem_result_29,
                   vinp2mem_result_30,
                   vinp2mem_result_31,
                   vinp2mem_result_32,
                   vinp2mem_result_33,
                   vinp2mem_result_34,
                   vinp2mem_result_35,
                   vinp2mem_result_36,
                   vinp2mem_result_37,
                   vinp2mem_result_38,
                   vinp2mem_result_39,
                   vinp2mem_result_40,
                   vinp2mem_result_41,
                   vinp2mem_result_42,
                   vinp2mem_result_43,
                   vinp2mem_result_44,
                   vinp2mem_result_45,
                   vinp2mem_result_46,
                   vinp2mem_result_47,
                   vinp2mem_result_48,
                   vinp2mem_result_49,
                   vinp2mem_result_50,
                   vinp2mem_result_51,
                   vinp2mem_result_52,
                   vinp2mem_result_53,
                   vinp2mem_result_54,
                   vinp2mem_result_55,
                   vinp2mem_result_56,
                   vinp2mem_result_57,
                   vinp2mem_result_58,
                   vinp2mem_result_59,
                   vinp2mem_result_60,
                   vinp2mem_result_61,
                   vinp2mem_result_62,
                   vinp2mem_result_63);
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_0;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_1;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_2;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_3;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_4;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_5;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_6;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_7;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_8;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_9;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_10;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_11;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_12;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_13;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_14;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_15;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_16;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_17;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_18;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_19;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_20;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_21;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_22;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_23;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_24;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_25;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_26;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_27;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_28;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_29;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_30;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_31;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_32;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_33;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_34;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_35;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_36;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_37;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_38;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_39;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_40;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_41;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_42;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_43;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_44;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_45;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_46;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_47;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_48;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_49;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_50;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_51;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_52;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_53;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_54;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_55;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_56;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_57;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_58;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_59;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_60;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_61;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_62;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_a_63;

    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_0;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_1;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_2;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_3;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_4;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_5;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_6;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_7;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_8;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_9;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_10;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_11;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_12;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_13;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_14;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_15;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_16;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_17;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_18;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_19;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_20;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_21;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_22;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_23;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_24;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_25;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_26;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_27;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_28;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_29;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_30;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_31;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_32;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_33;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_34;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_35;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_36;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_37;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_38;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_39;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_40;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_41;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_42;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_43;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_44;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_45;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_46;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_47;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_48;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_49;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_50;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_51;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_52;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_53;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_54;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_55;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_56;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_57;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_58;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_59;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_60;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_61;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_62;
    input       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     mem2vinp_b_63;

    input       [31:0]                          mem2vinp_size;

    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_0;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_1;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_2;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_3;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_4;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_5;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_6;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_7;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_8;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_9;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_10;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_11;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_12;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_13;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_14;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_15;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_16;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_17;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_18;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_19;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_20;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_21;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_22;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_23;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_24;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_25;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_26;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_27;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_28;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_29;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_30;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_31;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_32;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_33;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_34;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_35;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_36;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_37;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_38;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_39;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_40;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_41;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_42;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_43;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_44;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_45;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_46;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_47;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_48;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_49;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_50;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_51;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_52;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_53;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_54;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_55;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_56;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_57;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_58;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_59;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_60;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_61;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_62;
    output logic[`YTYDLA_mem2vinpA_LENGTH - 1:0]     vinp2mem_result_63;


    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_0;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_1;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_2;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_3;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_4;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_5;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_6;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_7;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_8;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_9;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_10;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_11;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_12;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_13;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_14;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_15;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_16;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_17;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_18;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_19;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_20;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_21;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_22;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_23;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_24;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_25;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_26;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_27;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_28;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_29;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_30;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_31;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_32;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_33;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_34;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_35;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_36;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_37;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_38;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_39;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_40;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_41;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_42;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_43;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_44;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_45;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_46;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_47;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_48;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_49;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_50;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_51;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_52;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_53;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_54;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_55;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_56;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_57;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_58;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_59;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_60;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_61;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_62;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_a_63;


    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_0;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_1;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_2;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_3;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_4;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_5;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_6;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_7;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_8;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_9;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_10;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_11;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_12;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_13;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_14;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_15;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_16;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_17;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_18;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_19;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_20;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_21;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_22;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_23;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_24;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_25;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_26;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_27;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_28;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_29;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_30;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_31;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_32;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_33;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_34;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_35;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_36;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_37;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_38;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_39;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_40;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_41;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_42;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_43;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_44;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_45;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_46;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_47;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_48;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_49;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_50;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_51;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_52;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_53;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_54;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_55;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_56;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_57;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_58;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_59;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_60;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_61;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_62;
    logic       [`YTYDLA_mem2vinpA_LENGTH - 1:0]     dat_b_63;



    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_0 <= 0;
        end
        if (mem2vinp_size > 0)begin
            dat_a_0 <= mem2vinp_a_0;
        end
        else begin
            dat_a_0 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_1 <= 0;
        end
        if (mem2vinp_size > 1)begin
            dat_a_1 <= mem2vinp_a_1;
        end
        else begin
            dat_a_1 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_2 <= 0;
        end
        if (mem2vinp_size > 2)begin
            dat_a_2 <= mem2vinp_a_2;
        end
        else begin
            dat_a_2 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_3 <= 0;
        end
        if (mem2vinp_size > 3)begin
            dat_a_3 <= mem2vinp_a_3;
        end
        else begin
            dat_a_3 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_4 <= 0;
        end
        if (mem2vinp_size > 4)begin
            dat_a_4 <= mem2vinp_a_4;
        end
        else begin
            dat_a_4 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_5 <= 0;
        end
        if (mem2vinp_size > 5)begin
            dat_a_5 <= mem2vinp_a_5;
        end
        else begin
            dat_a_5 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_6 <= 0;
        end
        if (mem2vinp_size > 6)begin
            dat_a_6 <= mem2vinp_a_6;
        end
        else begin
            dat_a_6 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_7 <= 0;
        end
        if (mem2vinp_size > 7)begin
            dat_a_7 <= mem2vinp_a_7;
        end
        else begin
            dat_a_7 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_8 <= 0;
        end
        if (mem2vinp_size > 8)begin
            dat_a_8 <= mem2vinp_a_8;
        end
        else begin
            dat_a_8 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_9 <= 0;
        end
        if (mem2vinp_size > 9)begin
            dat_a_9 <= mem2vinp_a_9;
        end
        else begin
            dat_a_9 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_10 <= 0;
        end
        if (mem2vinp_size > 10)begin
            dat_a_10 <= mem2vinp_a_10;
        end
        else begin
            dat_a_10 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_11 <= 0;
        end
        if (mem2vinp_size > 11)begin
            dat_a_11 <= mem2vinp_a_11;
        end
        else begin
            dat_a_11 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_12 <= 0;
        end
        if (mem2vinp_size > 12)begin
            dat_a_12 <= mem2vinp_a_12;
        end
        else begin
            dat_a_12 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_13 <= 0;
        end
        if (mem2vinp_size > 13)begin
            dat_a_13 <= mem2vinp_a_13;
        end
        else begin
            dat_a_13 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_14 <= 0;
        end
        if (mem2vinp_size > 14)begin
            dat_a_14 <= mem2vinp_a_14;
        end
        else begin
            dat_a_14 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_15 <= 0;
        end
        if (mem2vinp_size > 15)begin
            dat_a_15 <= mem2vinp_a_15;
        end
        else begin
            dat_a_15 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_16 <= 0;
        end
        if (mem2vinp_size > 16)begin
            dat_a_16 <= mem2vinp_a_16;
        end
        else begin
            dat_a_16 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_17 <= 0;
        end
        if (mem2vinp_size > 17)begin
            dat_a_17 <= mem2vinp_a_17;
        end
        else begin
            dat_a_17 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_18 <= 0;
        end
        if (mem2vinp_size > 18)begin
            dat_a_18 <= mem2vinp_a_18;
        end
        else begin
            dat_a_18 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_19 <= 0;
        end
        if (mem2vinp_size > 19)begin
            dat_a_19 <= mem2vinp_a_19;
        end
        else begin
            dat_a_19 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_20 <= 0;
        end
        if (mem2vinp_size > 20)begin
            dat_a_20 <= mem2vinp_a_20;
        end
        else begin
            dat_a_20 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_21 <= 0;
        end
        if (mem2vinp_size > 21)begin
            dat_a_21 <= mem2vinp_a_21;
        end
        else begin
            dat_a_21 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_22 <= 0;
        end
        if (mem2vinp_size > 22)begin
            dat_a_22 <= mem2vinp_a_22;
        end
        else begin
            dat_a_22 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_23 <= 0;
        end
        if (mem2vinp_size > 23)begin
            dat_a_23 <= mem2vinp_a_23;
        end
        else begin
            dat_a_23 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_24 <= 0;
        end
        if (mem2vinp_size > 24)begin
            dat_a_24 <= mem2vinp_a_24;
        end
        else begin
            dat_a_24 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_25 <= 0;
        end
        if (mem2vinp_size > 25)begin
            dat_a_25 <= mem2vinp_a_25;
        end
        else begin
            dat_a_25 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_26 <= 0;
        end
        if (mem2vinp_size > 26)begin
            dat_a_26 <= mem2vinp_a_26;
        end
        else begin
            dat_a_26 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_27 <= 0;
        end
        if (mem2vinp_size > 27)begin
            dat_a_27 <= mem2vinp_a_27;
        end
        else begin
            dat_a_27 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_28 <= 0;
        end
        if (mem2vinp_size > 28)begin
            dat_a_28 <= mem2vinp_a_28;
        end
        else begin
            dat_a_28 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_29 <= 0;
        end
        if (mem2vinp_size > 29)begin
            dat_a_29 <= mem2vinp_a_29;
        end
        else begin
            dat_a_29 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_30 <= 0;
        end
        if (mem2vinp_size > 30)begin
            dat_a_30 <= mem2vinp_a_30;
        end
        else begin
            dat_a_30 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_31 <= 0;
        end
        if (mem2vinp_size > 31)begin
            dat_a_31 <= mem2vinp_a_31;
        end
        else begin
            dat_a_31 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_32 <= 0;
        end
        if (mem2vinp_size > 32)begin
            dat_a_32 <= mem2vinp_a_32;
        end
        else begin
            dat_a_32 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_33 <= 0;
        end
        if (mem2vinp_size > 33)begin
            dat_a_33 <= mem2vinp_a_33;
        end
        else begin
            dat_a_33 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_34 <= 0;
        end
        if (mem2vinp_size > 34)begin
            dat_a_34 <= mem2vinp_a_34;
        end
        else begin
            dat_a_34 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_35 <= 0;
        end
        if (mem2vinp_size > 35)begin
            dat_a_35 <= mem2vinp_a_35;
        end
        else begin
            dat_a_35 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_36 <= 0;
        end
        if (mem2vinp_size > 36)begin
            dat_a_36 <= mem2vinp_a_36;
        end
        else begin
            dat_a_36 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_37 <= 0;
        end
        if (mem2vinp_size > 37)begin
            dat_a_37 <= mem2vinp_a_37;
        end
        else begin
            dat_a_37 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_38 <= 0;
        end
        if (mem2vinp_size > 38)begin
            dat_a_38 <= mem2vinp_a_38;
        end
        else begin
            dat_a_38 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_39 <= 0;
        end
        if (mem2vinp_size > 39)begin
            dat_a_39 <= mem2vinp_a_39;
        end
        else begin
            dat_a_39 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_40 <= 0;
        end
        if (mem2vinp_size > 40)begin
            dat_a_40 <= mem2vinp_a_40;
        end
        else begin
            dat_a_40 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_41 <= 0;
        end
        if (mem2vinp_size > 41)begin
            dat_a_41 <= mem2vinp_a_41;
        end
        else begin
            dat_a_41 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_42 <= 0;
        end
        if (mem2vinp_size > 42)begin
            dat_a_42 <= mem2vinp_a_42;
        end
        else begin
            dat_a_42 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_43 <= 0;
        end
        if (mem2vinp_size > 43)begin
            dat_a_43 <= mem2vinp_a_43;
        end
        else begin
            dat_a_43 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_44 <= 0;
        end
        if (mem2vinp_size > 44)begin
            dat_a_44 <= mem2vinp_a_44;
        end
        else begin
            dat_a_44 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_45 <= 0;
        end
        if (mem2vinp_size > 45)begin
            dat_a_45 <= mem2vinp_a_45;
        end
        else begin
            dat_a_45 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_46 <= 0;
        end
        if (mem2vinp_size > 46)begin
            dat_a_46 <= mem2vinp_a_46;
        end
        else begin
            dat_a_46 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_47 <= 0;
        end
        if (mem2vinp_size > 47)begin
            dat_a_47 <= mem2vinp_a_47;
        end
        else begin
            dat_a_47 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_48 <= 0;
        end
        if (mem2vinp_size > 48)begin
            dat_a_48 <= mem2vinp_a_48;
        end
        else begin
            dat_a_48 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_49 <= 0;
        end
        if (mem2vinp_size > 49)begin
            dat_a_49 <= mem2vinp_a_49;
        end
        else begin
            dat_a_49 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_50 <= 0;
        end
        if (mem2vinp_size > 50)begin
            dat_a_50 <= mem2vinp_a_50;
        end
        else begin
            dat_a_50 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_51 <= 0;
        end
        if (mem2vinp_size > 51)begin
            dat_a_51 <= mem2vinp_a_51;
        end
        else begin
            dat_a_51 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_52 <= 0;
        end
        if (mem2vinp_size > 52)begin
            dat_a_52 <= mem2vinp_a_52;
        end
        else begin
            dat_a_52 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_53 <= 0;
        end
        if (mem2vinp_size > 53)begin
            dat_a_53 <= mem2vinp_a_53;
        end
        else begin
            dat_a_53 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_54 <= 0;
        end
        if (mem2vinp_size > 54)begin
            dat_a_54 <= mem2vinp_a_54;
        end
        else begin
            dat_a_54 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_55 <= 0;
        end
        if (mem2vinp_size > 55)begin
            dat_a_55 <= mem2vinp_a_55;
        end
        else begin
            dat_a_55 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_56 <= 0;
        end
        if (mem2vinp_size > 56)begin
            dat_a_56 <= mem2vinp_a_56;
        end
        else begin
            dat_a_56 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_57 <= 0;
        end
        if (mem2vinp_size > 57)begin
            dat_a_57 <= mem2vinp_a_57;
        end
        else begin
            dat_a_57 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_58 <= 0;
        end
        if (mem2vinp_size > 58)begin
            dat_a_58 <= mem2vinp_a_58;
        end
        else begin
            dat_a_58 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_59 <= 0;
        end
        if (mem2vinp_size > 59)begin
            dat_a_59 <= mem2vinp_a_59;
        end
        else begin
            dat_a_59 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_60 <= 0;
        end
        if (mem2vinp_size > 60)begin
            dat_a_60 <= mem2vinp_a_60;
        end
        else begin
            dat_a_60 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_61 <= 0;
        end
        if (mem2vinp_size > 61)begin
            dat_a_61 <= mem2vinp_a_61;
        end
        else begin
            dat_a_61 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_62 <= 0;
        end
        if (mem2vinp_size > 62)begin
            dat_a_62 <= mem2vinp_a_62;
        end
        else begin
            dat_a_62 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_a_63 <= 0;
        end
        if (mem2vinp_size > 63)begin
            dat_a_63 <= mem2vinp_a_63;
        end
        else begin
            dat_a_63 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_0 <= 0;
        end
        if (mem2vinp_size > 0)begin
            dat_b_0 <= mem2vinp_b_0;
        end
        else begin
            dat_b_0 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_1 <= 0;
        end
        if (mem2vinp_size > 1)begin
            dat_b_1 <= mem2vinp_b_1;
        end
        else begin
            dat_b_1 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_2 <= 0;
        end
        if (mem2vinp_size > 2)begin
            dat_b_2 <= mem2vinp_b_2;
        end
        else begin
            dat_b_2 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_3 <= 0;
        end
        if (mem2vinp_size > 3)begin
            dat_b_3 <= mem2vinp_b_3;
        end
        else begin
            dat_b_3 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_4 <= 0;
        end
        if (mem2vinp_size > 4)begin
            dat_b_4 <= mem2vinp_b_4;
        end
        else begin
            dat_b_4 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_5 <= 0;
        end
        if (mem2vinp_size > 5)begin
            dat_b_5 <= mem2vinp_b_5;
        end
        else begin
            dat_b_5 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_6 <= 0;
        end
        if (mem2vinp_size > 6)begin
            dat_b_6 <= mem2vinp_b_6;
        end
        else begin
            dat_b_6 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_7 <= 0;
        end
        if (mem2vinp_size > 7)begin
            dat_b_7 <= mem2vinp_b_7;
        end
        else begin
            dat_b_7 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_8 <= 0;
        end
        if (mem2vinp_size > 8)begin
            dat_b_8 <= mem2vinp_b_8;
        end
        else begin
            dat_b_8 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_9 <= 0;
        end
        if (mem2vinp_size > 9)begin
            dat_b_9 <= mem2vinp_b_9;
        end
        else begin
            dat_b_9 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_10 <= 0;
        end
        if (mem2vinp_size > 10)begin
            dat_b_10 <= mem2vinp_b_10;
        end
        else begin
            dat_b_10 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_11 <= 0;
        end
        if (mem2vinp_size > 11)begin
            dat_b_11 <= mem2vinp_b_11;
        end
        else begin
            dat_b_11 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_12 <= 0;
        end
        if (mem2vinp_size > 12)begin
            dat_b_12 <= mem2vinp_b_12;
        end
        else begin
            dat_b_12 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_13 <= 0;
        end
        if (mem2vinp_size > 13)begin
            dat_b_13 <= mem2vinp_b_13;
        end
        else begin
            dat_b_13 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_14 <= 0;
        end
        if (mem2vinp_size > 14)begin
            dat_b_14 <= mem2vinp_b_14;
        end
        else begin
            dat_b_14 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_15 <= 0;
        end
        if (mem2vinp_size > 15)begin
            dat_b_15 <= mem2vinp_b_15;
        end
        else begin
            dat_b_15 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_16 <= 0;
        end
        if (mem2vinp_size > 16)begin
            dat_b_16 <= mem2vinp_b_16;
        end
        else begin
            dat_b_16 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_17 <= 0;
        end
        if (mem2vinp_size > 17)begin
            dat_b_17 <= mem2vinp_b_17;
        end
        else begin
            dat_b_17 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_18 <= 0;
        end
        if (mem2vinp_size > 18)begin
            dat_b_18 <= mem2vinp_b_18;
        end
        else begin
            dat_b_18 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_19 <= 0;
        end
        if (mem2vinp_size > 19)begin
            dat_b_19 <= mem2vinp_b_19;
        end
        else begin
            dat_b_19 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_20 <= 0;
        end
        if (mem2vinp_size > 20)begin
            dat_b_20 <= mem2vinp_b_20;
        end
        else begin
            dat_b_20 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_21 <= 0;
        end
        if (mem2vinp_size > 21)begin
            dat_b_21 <= mem2vinp_b_21;
        end
        else begin
            dat_b_21 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_22 <= 0;
        end
        if (mem2vinp_size > 22)begin
            dat_b_22 <= mem2vinp_b_22;
        end
        else begin
            dat_b_22 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_23 <= 0;
        end
        if (mem2vinp_size > 23)begin
            dat_b_23 <= mem2vinp_b_23;
        end
        else begin
            dat_b_23 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_24 <= 0;
        end
        if (mem2vinp_size > 24)begin
            dat_b_24 <= mem2vinp_b_24;
        end
        else begin
            dat_b_24 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_25 <= 0;
        end
        if (mem2vinp_size > 25)begin
            dat_b_25 <= mem2vinp_b_25;
        end
        else begin
            dat_b_25 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_26 <= 0;
        end
        if (mem2vinp_size > 26)begin
            dat_b_26 <= mem2vinp_b_26;
        end
        else begin
            dat_b_26 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_27 <= 0;
        end
        if (mem2vinp_size > 27)begin
            dat_b_27 <= mem2vinp_b_27;
        end
        else begin
            dat_b_27 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_28 <= 0;
        end
        if (mem2vinp_size > 28)begin
            dat_b_28 <= mem2vinp_b_28;
        end
        else begin
            dat_b_28 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_29 <= 0;
        end
        if (mem2vinp_size > 29)begin
            dat_b_29 <= mem2vinp_b_29;
        end
        else begin
            dat_b_29 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_30 <= 0;
        end
        if (mem2vinp_size > 30)begin
            dat_b_30 <= mem2vinp_b_30;
        end
        else begin
            dat_b_30 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_31 <= 0;
        end
        if (mem2vinp_size > 31)begin
            dat_b_31 <= mem2vinp_b_31;
        end
        else begin
            dat_b_31 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_32 <= 0;
        end
        if (mem2vinp_size > 32)begin
            dat_b_32 <= mem2vinp_b_32;
        end
        else begin
            dat_b_32 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_33 <= 0;
        end
        if (mem2vinp_size > 33)begin
            dat_b_33 <= mem2vinp_b_33;
        end
        else begin
            dat_b_33 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_34 <= 0;
        end
        if (mem2vinp_size > 34)begin
            dat_b_34 <= mem2vinp_b_34;
        end
        else begin
            dat_b_34 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_35 <= 0;
        end
        if (mem2vinp_size > 35)begin
            dat_b_35 <= mem2vinp_b_35;
        end
        else begin
            dat_b_35 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_36 <= 0;
        end
        if (mem2vinp_size > 36)begin
            dat_b_36 <= mem2vinp_b_36;
        end
        else begin
            dat_b_36 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_37 <= 0;
        end
        if (mem2vinp_size > 37)begin
            dat_b_37 <= mem2vinp_b_37;
        end
        else begin
            dat_b_37 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_38 <= 0;
        end
        if (mem2vinp_size > 38)begin
            dat_b_38 <= mem2vinp_b_38;
        end
        else begin
            dat_b_38 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_39 <= 0;
        end
        if (mem2vinp_size > 39)begin
            dat_b_39 <= mem2vinp_b_39;
        end
        else begin
            dat_b_39 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_40 <= 0;
        end
        if (mem2vinp_size > 40)begin
            dat_b_40 <= mem2vinp_b_40;
        end
        else begin
            dat_b_40 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_41 <= 0;
        end
        if (mem2vinp_size > 41)begin
            dat_b_41 <= mem2vinp_b_41;
        end
        else begin
            dat_b_41 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_42 <= 0;
        end
        if (mem2vinp_size > 42)begin
            dat_b_42 <= mem2vinp_b_42;
        end
        else begin
            dat_b_42 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_43 <= 0;
        end
        if (mem2vinp_size > 43)begin
            dat_b_43 <= mem2vinp_b_43;
        end
        else begin
            dat_b_43 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_44 <= 0;
        end
        if (mem2vinp_size > 44)begin
            dat_b_44 <= mem2vinp_b_44;
        end
        else begin
            dat_b_44 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_45 <= 0;
        end
        if (mem2vinp_size > 45)begin
            dat_b_45 <= mem2vinp_b_45;
        end
        else begin
            dat_b_45 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_46 <= 0;
        end
        if (mem2vinp_size > 46)begin
            dat_b_46 <= mem2vinp_b_46;
        end
        else begin
            dat_b_46 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_47 <= 0;
        end
        if (mem2vinp_size > 47)begin
            dat_b_47 <= mem2vinp_b_47;
        end
        else begin
            dat_b_47 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_48 <= 0;
        end
        if (mem2vinp_size > 48)begin
            dat_b_48 <= mem2vinp_b_48;
        end
        else begin
            dat_b_48 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_49 <= 0;
        end
        if (mem2vinp_size > 49)begin
            dat_b_49 <= mem2vinp_b_49;
        end
        else begin
            dat_b_49 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_50 <= 0;
        end
        if (mem2vinp_size > 50)begin
            dat_b_50 <= mem2vinp_b_50;
        end
        else begin
            dat_b_50 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_51 <= 0;
        end
        if (mem2vinp_size > 51)begin
            dat_b_51 <= mem2vinp_b_51;
        end
        else begin
            dat_b_51 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_52 <= 0;
        end
        if (mem2vinp_size > 52)begin
            dat_b_52 <= mem2vinp_b_52;
        end
        else begin
            dat_b_52 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_53 <= 0;
        end
        if (mem2vinp_size > 53)begin
            dat_b_53 <= mem2vinp_b_53;
        end
        else begin
            dat_b_53 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_54 <= 0;
        end
        if (mem2vinp_size > 54)begin
            dat_b_54 <= mem2vinp_b_54;
        end
        else begin
            dat_b_54 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_55 <= 0;
        end
        if (mem2vinp_size > 55)begin
            dat_b_55 <= mem2vinp_b_55;
        end
        else begin
            dat_b_55 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_56 <= 0;
        end
        if (mem2vinp_size > 56)begin
            dat_b_56 <= mem2vinp_b_56;
        end
        else begin
            dat_b_56 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_57 <= 0;
        end
        if (mem2vinp_size > 57)begin
            dat_b_57 <= mem2vinp_b_57;
        end
        else begin
            dat_b_57 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_58 <= 0;
        end
        if (mem2vinp_size > 58)begin
            dat_b_58 <= mem2vinp_b_58;
        end
        else begin
            dat_b_58 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_59 <= 0;
        end
        if (mem2vinp_size > 59)begin
            dat_b_59 <= mem2vinp_b_59;
        end
        else begin
            dat_b_59 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_60 <= 0;
        end
        if (mem2vinp_size > 60)begin
            dat_b_60 <= mem2vinp_b_60;
        end
        else begin
            dat_b_60 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_61 <= 0;
        end
        if (mem2vinp_size > 61)begin
            dat_b_61 <= mem2vinp_b_61;
        end
        else begin
            dat_b_61 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_62 <= 0;
        end
        if (mem2vinp_size > 62)begin
            dat_b_62 <= mem2vinp_b_62;
        end
        else begin
            dat_b_62 <= 0;
        end
    end

    always_ff @(posedge ytydla_core_clk or negedge ytydla_core_rst_n)begin
        if (~ytydla_core_rst_n)begin
            dat_b_63 <= 0;
        end
        if (mem2vinp_size > 63)begin
            dat_b_63 <= mem2vinp_b_63;
        end
        else begin
            dat_b_63 <= 0;
        end
    end

    ytydla_cmac_mul    mul_0(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_0),
                          .weight (dat_b_0),
                          .result (vinp2mem_result_0));
    ytydla_cmac_mul    mul_1(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_1),
                          .weight (dat_b_1),
                          .result (vinp2mem_result_1));
    ytydla_cmac_mul    mul_2(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_2),
                          .weight (dat_b_2),
                          .result (vinp2mem_result_2));
    ytydla_cmac_mul    mul_3(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_3),
                          .weight (dat_b_3),
                          .result (vinp2mem_result_3));
    ytydla_cmac_mul    mul_4(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_4),
                          .weight (dat_b_4),
                          .result (vinp2mem_result_4));
    ytydla_cmac_mul    mul_5(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_5),
                          .weight (dat_b_5),
                          .result (vinp2mem_result_5));
    ytydla_cmac_mul    mul_6(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_6),
                          .weight (dat_b_6),
                          .result (vinp2mem_result_6));
    ytydla_cmac_mul    mul_7(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_7),
                          .weight (dat_b_7),
                          .result (vinp2mem_result_7));
    ytydla_cmac_mul    mul_8(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_8),
                          .weight (dat_b_8),
                          .result (vinp2mem_result_8));
    ytydla_cmac_mul    mul_9(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_9),
                          .weight (dat_b_9),
                          .result (vinp2mem_result_9));
    ytydla_cmac_mul    mul_10(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_10),
                          .weight (dat_b_10),
                          .result (vinp2mem_result_10));
    ytydla_cmac_mul    mul_11(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_11),
                          .weight (dat_b_11),
                          .result (vinp2mem_result_11));
    ytydla_cmac_mul    mul_12(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_12),
                          .weight (dat_b_12),
                          .result (vinp2mem_result_12));
    ytydla_cmac_mul    mul_13(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_13),
                          .weight (dat_b_13),
                          .result (vinp2mem_result_13));
    ytydla_cmac_mul    mul_14(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_14),
                          .weight (dat_b_14),
                          .result (vinp2mem_result_14));
    ytydla_cmac_mul    mul_15(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_15),
                          .weight (dat_b_15),
                          .result (vinp2mem_result_15));
    ytydla_cmac_mul    mul_16(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_16),
                          .weight (dat_b_16),
                          .result (vinp2mem_result_16));
    ytydla_cmac_mul    mul_17(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_17),
                          .weight (dat_b_17),
                          .result (vinp2mem_result_17));
    ytydla_cmac_mul    mul_18(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_18),
                          .weight (dat_b_18),
                          .result (vinp2mem_result_18));
    ytydla_cmac_mul    mul_19(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_19),
                          .weight (dat_b_19),
                          .result (vinp2mem_result_19));
    ytydla_cmac_mul    mul_20(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_20),
                          .weight (dat_b_20),
                          .result (vinp2mem_result_20));
    ytydla_cmac_mul    mul_21(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_21),
                          .weight (dat_b_21),
                          .result (vinp2mem_result_21));
    ytydla_cmac_mul    mul_22(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_22),
                          .weight (dat_b_22),
                          .result (vinp2mem_result_22));
    ytydla_cmac_mul    mul_23(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_23),
                          .weight (dat_b_23),
                          .result (vinp2mem_result_23));
    ytydla_cmac_mul    mul_24(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_24),
                          .weight (dat_b_24),
                          .result (vinp2mem_result_24));
    ytydla_cmac_mul    mul_25(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_25),
                          .weight (dat_b_25),
                          .result (vinp2mem_result_25));
    ytydla_cmac_mul    mul_26(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_26),
                          .weight (dat_b_26),
                          .result (vinp2mem_result_26));
    ytydla_cmac_mul    mul_27(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_27),
                          .weight (dat_b_27),
                          .result (vinp2mem_result_27));
    ytydla_cmac_mul    mul_28(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_28),
                          .weight (dat_b_28),
                          .result (vinp2mem_result_28));
    ytydla_cmac_mul    mul_29(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_29),
                          .weight (dat_b_29),
                          .result (vinp2mem_result_29));
    ytydla_cmac_mul    mul_30(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_30),
                          .weight (dat_b_30),
                          .result (vinp2mem_result_30));
    ytydla_cmac_mul    mul_31(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_31),
                          .weight (dat_b_31),
                          .result (vinp2mem_result_31));
    ytydla_cmac_mul    mul_32(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_32),
                          .weight (dat_b_32),
                          .result (vinp2mem_result_32));
    ytydla_cmac_mul    mul_33(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_33),
                          .weight (dat_b_33),
                          .result (vinp2mem_result_33));
    ytydla_cmac_mul    mul_34(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_34),
                          .weight (dat_b_34),
                          .result (vinp2mem_result_34));
    ytydla_cmac_mul    mul_35(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_35),
                          .weight (dat_b_35),
                          .result (vinp2mem_result_35));
    ytydla_cmac_mul    mul_36(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_36),
                          .weight (dat_b_36),
                          .result (vinp2mem_result_36));
    ytydla_cmac_mul    mul_37(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_37),
                          .weight (dat_b_37),
                          .result (vinp2mem_result_37));
    ytydla_cmac_mul    mul_38(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_38),
                          .weight (dat_b_38),
                          .result (vinp2mem_result_38));
    ytydla_cmac_mul    mul_39(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_39),
                          .weight (dat_b_39),
                          .result (vinp2mem_result_39));
    ytydla_cmac_mul    mul_40(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_40),
                          .weight (dat_b_40),
                          .result (vinp2mem_result_40));
    ytydla_cmac_mul    mul_41(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_41),
                          .weight (dat_b_41),
                          .result (vinp2mem_result_41));
    ytydla_cmac_mul    mul_42(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_42),
                          .weight (dat_b_42),
                          .result (vinp2mem_result_42));
    ytydla_cmac_mul    mul_43(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_43),
                          .weight (dat_b_43),
                          .result (vinp2mem_result_43));
    ytydla_cmac_mul    mul_44(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_44),
                          .weight (dat_b_44),
                          .result (vinp2mem_result_44));
    ytydla_cmac_mul    mul_45(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_45),
                          .weight (dat_b_45),
                          .result (vinp2mem_result_45));
    ytydla_cmac_mul    mul_46(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_46),
                          .weight (dat_b_46),
                          .result (vinp2mem_result_46));
    ytydla_cmac_mul    mul_47(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_47),
                          .weight (dat_b_47),
                          .result (vinp2mem_result_47));
    ytydla_cmac_mul    mul_48(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_48),
                          .weight (dat_b_48),
                          .result (vinp2mem_result_48));
    ytydla_cmac_mul    mul_49(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_49),
                          .weight (dat_b_49),
                          .result (vinp2mem_result_49));
    ytydla_cmac_mul    mul_50(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_50),
                          .weight (dat_b_50),
                          .result (vinp2mem_result_50));
    ytydla_cmac_mul    mul_51(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_51),
                          .weight (dat_b_51),
                          .result (vinp2mem_result_51));
    ytydla_cmac_mul    mul_52(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_52),
                          .weight (dat_b_52),
                          .result (vinp2mem_result_52));
    ytydla_cmac_mul    mul_53(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_53),
                          .weight (dat_b_53),
                          .result (vinp2mem_result_53));
    ytydla_cmac_mul    mul_54(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_54),
                          .weight (dat_b_54),
                          .result (vinp2mem_result_54));
    ytydla_cmac_mul    mul_55(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_55),
                          .weight (dat_b_55),
                          .result (vinp2mem_result_55));
    ytydla_cmac_mul    mul_56(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_56),
                          .weight (dat_b_56),
                          .result (vinp2mem_result_56));
    ytydla_cmac_mul    mul_57(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_57),
                          .weight (dat_b_57),
                          .result (vinp2mem_result_57));
    ytydla_cmac_mul    mul_58(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_58),
                          .weight (dat_b_58),
                          .result (vinp2mem_result_58));
    ytydla_cmac_mul    mul_59(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_59),
                          .weight (dat_b_59),
                          .result (vinp2mem_result_59));
    ytydla_cmac_mul    mul_60(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_60),
                          .weight (dat_b_60),
                          .result (vinp2mem_result_60));
    ytydla_cmac_mul    mul_61(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_61),
                          .weight (dat_b_61),
                          .result (vinp2mem_result_61));
    ytydla_cmac_mul    mul_62(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_62),
                          .weight (dat_b_62),
                          .result (vinp2mem_result_62));
    ytydla_cmac_mul    mul_63(.clk    (ytydla_core_clk),
                          .rst_n  (ytydla_core_rst_n),
                          .data   (dat_a_63),
                          .weight (dat_b_63),
                          .result (vinp2mem_result_63));

endmodule
