﻿//ytydla.sv


module ytydla_tb;
    integer i;
    logic   ytydla_core_clk;
    logic   ytydla_core_rst_n;
    logic [7:0] memory[0:65535];
    logic [31:0] data_size = 28;
    logic [31:0] weight_size = 5;
    $readmemh("data/memory.lists", memory);

    initial begin
        ytydla_core_clk = 0;
        ytydla_core_rst_n = 0;
        #1 ytydla_core_rst_n = 1;
        for (i = 0; i < 100; i = i + 1)begin
            #1 ytydla_core_clk = ~ytydla_core_clk;
        end
    ytydla_conv2d conv_0(
        .ytydla_core_clk    ytydla_core_clk,
        .ytydla_core_rst_n  ytydla_core_rst_n,
        .ls2cmac_dat0       {memory[3], memory[2], memory[1], memory[0]},
        .ls2cmac_dat1       {memory[7], memory[6], memory[5], memory[4]},
        .ls2cmac_dat2       {memory[11], memory[10], memory[9], memory[8]},
        .ls2cmac_dat3       {memory[15], memory[14], memory[13], memory[12]},
        .ls2cmac_dat4       {memory[19], memory[18], memory[17], memory[16]},
        .ls2cmac_dat5       {memory[23], memory[22], memory[21], memory[20]},
        .ls2cmac_dat6       {memory[27], memory[26], memory[25], memory[24]},
        .ls2cmac_dat7       {memory[31], memory[30], memory[29], memory[28]},
        .ls2cmac_dat8       {memory[35], memory[34], memory[33], memory[32]},
        .ls2cmac_dat9       {memory[39], memory[38], memory[37], memory[36]},
        .ls2cmac_dat10       {memory[43], memory[42], memory[41], memory[40]},
        .ls2cmac_dat11       {memory[47], memory[46], memory[45], memory[44]},
        .ls2cmac_dat12       {memory[51], memory[50], memory[49], memory[48]},
        .ls2cmac_dat13       {memory[55], memory[54], memory[53], memory[52]},
        .ls2cmac_dat14       {memory[59], memory[58], memory[57], memory[56]},
        .ls2cmac_dat15       {memory[63], memory[62], memory[61], memory[60]},
        .ls2cmac_dat16       {memory[67], memory[66], memory[65], memory[64]},
        .ls2cmac_dat17       {memory[71], memory[70], memory[69], memory[68]},
        .ls2cmac_dat18       {memory[75], memory[74], memory[73], memory[72]},
        .ls2cmac_dat19       {memory[79], memory[78], memory[77], memory[76]},
        .ls2cmac_dat20       {memory[83], memory[82], memory[81], memory[80]},
        .ls2cmac_dat21       {memory[87], memory[86], memory[85], memory[84]},
        .ls2cmac_dat22       {memory[91], memory[90], memory[89], memory[88]},
        .ls2cmac_dat23       {memory[95], memory[94], memory[93], memory[92]},
        .ls2cmac_dat24       {memory[99], memory[98], memory[97], memory[96]},
        .ls2cmac_dat25       {memory[103], memory[102], memory[101], memory[100]},
        .ls2cmac_dat26       {memory[107], memory[106], memory[105], memory[104]},
        .ls2cmac_dat27       {memory[111], memory[110], memory[109], memory[108]},
        .ls2cmac_dat28       {memory[115], memory[114], memory[113], memory[112]},
        .ls2cmac_dat29       {memory[119], memory[118], memory[117], memory[116]},
        .ls2cmac_dat30       {memory[123], memory[122], memory[121], memory[120]},
        .ls2cmac_dat31       {memory[127], memory[126], memory[125], memory[124]},
        .ls2cmac_dat32       {memory[131], memory[130], memory[129], memory[128]},
        .ls2cmac_dat33       {memory[135], memory[134], memory[133], memory[132]},
        .ls2cmac_dat34       {memory[139], memory[138], memory[137], memory[136]},
        .ls2cmac_dat35       {memory[143], memory[142], memory[141], memory[140]},
        .ls2cmac_dat36       {memory[147], memory[146], memory[145], memory[144]},
        .ls2cmac_dat37       {memory[151], memory[150], memory[149], memory[148]},
        .ls2cmac_dat38       {memory[155], memory[154], memory[153], memory[152]},
        .ls2cmac_dat39       {memory[159], memory[158], memory[157], memory[156]},
        .ls2cmac_dat40       {memory[163], memory[162], memory[161], memory[160]},
        .ls2cmac_dat41       {memory[167], memory[166], memory[165], memory[164]},
        .ls2cmac_dat42       {memory[171], memory[170], memory[169], memory[168]},
        .ls2cmac_dat43       {memory[175], memory[174], memory[173], memory[172]},
        .ls2cmac_dat44       {memory[179], memory[178], memory[177], memory[176]},
        .ls2cmac_dat45       {memory[183], memory[182], memory[181], memory[180]},
        .ls2cmac_dat46       {memory[187], memory[186], memory[185], memory[184]},
        .ls2cmac_dat47       {memory[191], memory[190], memory[189], memory[188]},
        .ls2cmac_dat48       {memory[195], memory[194], memory[193], memory[192]},
        .ls2cmac_dat49       {memory[199], memory[198], memory[197], memory[196]},
        .ls2cmac_dat50       {memory[203], memory[202], memory[201], memory[200]},
        .ls2cmac_dat51       {memory[207], memory[206], memory[205], memory[204]},
        .ls2cmac_dat52       {memory[211], memory[210], memory[209], memory[208]},
        .ls2cmac_dat53       {memory[215], memory[214], memory[213], memory[212]},
        .ls2cmac_dat54       {memory[219], memory[218], memory[217], memory[216]},
        .ls2cmac_dat55       {memory[223], memory[222], memory[221], memory[220]},
        .ls2cmac_dat56       {memory[227], memory[226], memory[225], memory[224]},
        .ls2cmac_dat57       {memory[231], memory[230], memory[229], memory[228]},
        .ls2cmac_dat58       {memory[235], memory[234], memory[233], memory[232]},
        .ls2cmac_dat59       {memory[239], memory[238], memory[237], memory[236]},
        .ls2cmac_dat60       {memory[243], memory[242], memory[241], memory[240]},
        .ls2cmac_dat61       {memory[247], memory[246], memory[245], memory[244]},
        .ls2cmac_dat62       {memory[251], memory[250], memory[249], memory[248]},
        .ls2cmac_dat63       {memory[255], memory[254], memory[253], memory[252]},
        .ls2cmac_dat64       {memory[259], memory[258], memory[257], memory[256]},
        .ls2cmac_dat65       {memory[263], memory[262], memory[261], memory[260]},
        .ls2cmac_dat66       {memory[267], memory[266], memory[265], memory[264]},
        .ls2cmac_dat67       {memory[271], memory[270], memory[269], memory[268]},
        .ls2cmac_dat68       {memory[275], memory[274], memory[273], memory[272]},
        .ls2cmac_dat69       {memory[279], memory[278], memory[277], memory[276]},
        .ls2cmac_dat70       {memory[283], memory[282], memory[281], memory[280]},
        .ls2cmac_dat71       {memory[287], memory[286], memory[285], memory[284]},
        .ls2cmac_dat72       {memory[291], memory[290], memory[289], memory[288]},
        .ls2cmac_dat73       {memory[295], memory[294], memory[293], memory[292]},
        .ls2cmac_dat74       {memory[299], memory[298], memory[297], memory[296]},
        .ls2cmac_dat75       {memory[303], memory[302], memory[301], memory[300]},
        .ls2cmac_dat76       {memory[307], memory[306], memory[305], memory[304]},
        .ls2cmac_dat77       {memory[311], memory[310], memory[309], memory[308]},
        .ls2cmac_dat78       {memory[315], memory[314], memory[313], memory[312]},
        .ls2cmac_dat79       {memory[319], memory[318], memory[317], memory[316]},
        .ls2cmac_dat80       {memory[323], memory[322], memory[321], memory[320]},
        .ls2cmac_dat81       {memory[327], memory[326], memory[325], memory[324]},
        .ls2cmac_dat82       {memory[331], memory[330], memory[329], memory[328]},
        .ls2cmac_dat83       {memory[335], memory[334], memory[333], memory[332]},
        .ls2cmac_dat84       {memory[339], memory[338], memory[337], memory[336]},
        .ls2cmac_dat85       {memory[343], memory[342], memory[341], memory[340]},
        .ls2cmac_dat86       {memory[347], memory[346], memory[345], memory[344]},
        .ls2cmac_dat87       {memory[351], memory[350], memory[349], memory[348]},
        .ls2cmac_dat88       {memory[355], memory[354], memory[353], memory[352]},
        .ls2cmac_dat89       {memory[359], memory[358], memory[357], memory[356]},
        .ls2cmac_dat90       {memory[363], memory[362], memory[361], memory[360]},
        .ls2cmac_dat91       {memory[367], memory[366], memory[365], memory[364]},
        .ls2cmac_dat92       {memory[371], memory[370], memory[369], memory[368]},
        .ls2cmac_dat93       {memory[375], memory[374], memory[373], memory[372]},
        .ls2cmac_dat94       {memory[379], memory[378], memory[377], memory[376]},
        .ls2cmac_dat95       {memory[383], memory[382], memory[381], memory[380]},
        .ls2cmac_dat96       {memory[387], memory[386], memory[385], memory[384]},
        .ls2cmac_dat97       {memory[391], memory[390], memory[389], memory[388]},
        .ls2cmac_dat98       {memory[395], memory[394], memory[393], memory[392]},
        .ls2cmac_dat99       {memory[399], memory[398], memory[397], memory[396]},
        .ls2cmac_dat100       {memory[403], memory[402], memory[401], memory[400]},
        .ls2cmac_dat101       {memory[407], memory[406], memory[405], memory[404]},
        .ls2cmac_dat102       {memory[411], memory[410], memory[409], memory[408]},
        .ls2cmac_dat103       {memory[415], memory[414], memory[413], memory[412]},
        .ls2cmac_dat104       {memory[419], memory[418], memory[417], memory[416]},
        .ls2cmac_dat105       {memory[423], memory[422], memory[421], memory[420]},
        .ls2cmac_dat106       {memory[427], memory[426], memory[425], memory[424]},
        .ls2cmac_dat107       {memory[431], memory[430], memory[429], memory[428]},
        .ls2cmac_dat108       {memory[435], memory[434], memory[433], memory[432]},
        .ls2cmac_dat109       {memory[439], memory[438], memory[437], memory[436]},
        .ls2cmac_dat110       {memory[443], memory[442], memory[441], memory[440]},
        .ls2cmac_dat111       {memory[447], memory[446], memory[445], memory[444]},
        .ls2cmac_dat112       {memory[451], memory[450], memory[449], memory[448]},
        .ls2cmac_dat113       {memory[455], memory[454], memory[453], memory[452]},
        .ls2cmac_dat114       {memory[459], memory[458], memory[457], memory[456]},
        .ls2cmac_dat115       {memory[463], memory[462], memory[461], memory[460]},
        .ls2cmac_dat116       {memory[467], memory[466], memory[465], memory[464]},
        .ls2cmac_dat117       {memory[471], memory[470], memory[469], memory[468]},
        .ls2cmac_dat118       {memory[475], memory[474], memory[473], memory[472]},
        .ls2cmac_dat119       {memory[479], memory[478], memory[477], memory[476]},
        .ls2cmac_dat120       {memory[483], memory[482], memory[481], memory[480]},
        .ls2cmac_dat121       {memory[487], memory[486], memory[485], memory[484]},
        .ls2cmac_dat122       {memory[491], memory[490], memory[489], memory[488]},
        .ls2cmac_dat123       {memory[495], memory[494], memory[493], memory[492]},
        .ls2cmac_dat124       {memory[499], memory[498], memory[497], memory[496]},
        .ls2cmac_dat125       {memory[503], memory[502], memory[501], memory[500]},
        .ls2cmac_dat126       {memory[507], memory[506], memory[505], memory[504]},
        .ls2cmac_dat127       {memory[511], memory[510], memory[509], memory[508]},
        .ls2cmac_dat128       {memory[515], memory[514], memory[513], memory[512]},
        .ls2cmac_dat129       {memory[519], memory[518], memory[517], memory[516]},
        .ls2cmac_dat130       {memory[523], memory[522], memory[521], memory[520]},
        .ls2cmac_dat131       {memory[527], memory[526], memory[525], memory[524]},
        .ls2cmac_dat132       {memory[531], memory[530], memory[529], memory[528]},
        .ls2cmac_dat133       {memory[535], memory[534], memory[533], memory[532]},
        .ls2cmac_dat134       {memory[539], memory[538], memory[537], memory[536]},
        .ls2cmac_dat135       {memory[543], memory[542], memory[541], memory[540]},
        .ls2cmac_dat136       {memory[547], memory[546], memory[545], memory[544]},
        .ls2cmac_dat137       {memory[551], memory[550], memory[549], memory[548]},
        .ls2cmac_dat138       {memory[555], memory[554], memory[553], memory[552]},
        .ls2cmac_dat139       {memory[559], memory[558], memory[557], memory[556]},
        .ls2cmac_dat140       {memory[563], memory[562], memory[561], memory[560]},
        .ls2cmac_dat141       {memory[567], memory[566], memory[565], memory[564]},
        .ls2cmac_dat142       {memory[571], memory[570], memory[569], memory[568]},
        .ls2cmac_dat143       {memory[575], memory[574], memory[573], memory[572]},
        .ls2cmac_dat144       {memory[579], memory[578], memory[577], memory[576]},
        .ls2cmac_dat145       {memory[583], memory[582], memory[581], memory[580]},
        .ls2cmac_dat146       {memory[587], memory[586], memory[585], memory[584]},
        .ls2cmac_dat147       {memory[591], memory[590], memory[589], memory[588]},
        .ls2cmac_dat148       {memory[595], memory[594], memory[593], memory[592]},
        .ls2cmac_dat149       {memory[599], memory[598], memory[597], memory[596]},
        .ls2cmac_dat150       {memory[603], memory[602], memory[601], memory[600]},
        .ls2cmac_dat151       {memory[607], memory[606], memory[605], memory[604]},
        .ls2cmac_dat152       {memory[611], memory[610], memory[609], memory[608]},
        .ls2cmac_dat153       {memory[615], memory[614], memory[613], memory[612]},
        .ls2cmac_dat154       {memory[619], memory[618], memory[617], memory[616]},
        .ls2cmac_dat155       {memory[623], memory[622], memory[621], memory[620]},
        .ls2cmac_dat156       {memory[627], memory[626], memory[625], memory[624]},
        .ls2cmac_dat157       {memory[631], memory[630], memory[629], memory[628]},
        .ls2cmac_dat158       {memory[635], memory[634], memory[633], memory[632]},
        .ls2cmac_dat159       {memory[639], memory[638], memory[637], memory[636]},
        .ls2cmac_dat160       {memory[643], memory[642], memory[641], memory[640]},
        .ls2cmac_dat161       {memory[647], memory[646], memory[645], memory[644]},
        .ls2cmac_dat162       {memory[651], memory[650], memory[649], memory[648]},
        .ls2cmac_dat163       {memory[655], memory[654], memory[653], memory[652]},
        .ls2cmac_dat164       {memory[659], memory[658], memory[657], memory[656]},
        .ls2cmac_dat165       {memory[663], memory[662], memory[661], memory[660]},
        .ls2cmac_dat166       {memory[667], memory[666], memory[665], memory[664]},
        .ls2cmac_dat167       {memory[671], memory[670], memory[669], memory[668]},
        .ls2cmac_dat168       {memory[675], memory[674], memory[673], memory[672]},
        .ls2cmac_dat169       {memory[679], memory[678], memory[677], memory[676]},
        .ls2cmac_dat170       {memory[683], memory[682], memory[681], memory[680]},
        .ls2cmac_dat171       {memory[687], memory[686], memory[685], memory[684]},
        .ls2cmac_dat172       {memory[691], memory[690], memory[689], memory[688]},
        .ls2cmac_dat173       {memory[695], memory[694], memory[693], memory[692]},
        .ls2cmac_dat174       {memory[699], memory[698], memory[697], memory[696]},
        .ls2cmac_dat175       {memory[703], memory[702], memory[701], memory[700]},
        .ls2cmac_dat176       {memory[707], memory[706], memory[705], memory[704]},
        .ls2cmac_dat177       {memory[711], memory[710], memory[709], memory[708]},
        .ls2cmac_dat178       {memory[715], memory[714], memory[713], memory[712]},
        .ls2cmac_dat179       {memory[719], memory[718], memory[717], memory[716]},
        .ls2cmac_dat180       {memory[723], memory[722], memory[721], memory[720]},
        .ls2cmac_dat181       {memory[727], memory[726], memory[725], memory[724]},
        .ls2cmac_dat182       {memory[731], memory[730], memory[729], memory[728]},
        .ls2cmac_dat183       {memory[735], memory[734], memory[733], memory[732]},
        .ls2cmac_dat184       {memory[739], memory[738], memory[737], memory[736]},
        .ls2cmac_dat185       {memory[743], memory[742], memory[741], memory[740]},
        .ls2cmac_dat186       {memory[747], memory[746], memory[745], memory[744]},
        .ls2cmac_dat187       {memory[751], memory[750], memory[749], memory[748]},
        .ls2cmac_dat188       {memory[755], memory[754], memory[753], memory[752]},
        .ls2cmac_dat189       {memory[759], memory[758], memory[757], memory[756]},
        .ls2cmac_dat190       {memory[763], memory[762], memory[761], memory[760]},
        .ls2cmac_dat191       {memory[767], memory[766], memory[765], memory[764]},
        .ls2cmac_dat192       {memory[771], memory[770], memory[769], memory[768]},
        .ls2cmac_dat193       {memory[775], memory[774], memory[773], memory[772]},
        .ls2cmac_dat194       {memory[779], memory[778], memory[777], memory[776]},
        .ls2cmac_dat195       {memory[783], memory[782], memory[781], memory[780]},
        .ls2cmac_dat196       {memory[787], memory[786], memory[785], memory[784]},
        .ls2cmac_dat197       {memory[791], memory[790], memory[789], memory[788]},
        .ls2cmac_dat198       {memory[795], memory[794], memory[793], memory[792]},
        .ls2cmac_dat199       {memory[799], memory[798], memory[797], memory[796]},
        .ls2cmac_dat200       {memory[803], memory[802], memory[801], memory[800]},
        .ls2cmac_dat201       {memory[807], memory[806], memory[805], memory[804]},
        .ls2cmac_dat202       {memory[811], memory[810], memory[809], memory[808]},
        .ls2cmac_dat203       {memory[815], memory[814], memory[813], memory[812]},
        .ls2cmac_dat204       {memory[819], memory[818], memory[817], memory[816]},
        .ls2cmac_dat205       {memory[823], memory[822], memory[821], memory[820]},
        .ls2cmac_dat206       {memory[827], memory[826], memory[825], memory[824]},
        .ls2cmac_dat207       {memory[831], memory[830], memory[829], memory[828]},
        .ls2cmac_dat208       {memory[835], memory[834], memory[833], memory[832]},
        .ls2cmac_dat209       {memory[839], memory[838], memory[837], memory[836]},
        .ls2cmac_dat210       {memory[843], memory[842], memory[841], memory[840]},
        .ls2cmac_dat211       {memory[847], memory[846], memory[845], memory[844]},
        .ls2cmac_dat212       {memory[851], memory[850], memory[849], memory[848]},
        .ls2cmac_dat213       {memory[855], memory[854], memory[853], memory[852]},
        .ls2cmac_dat214       {memory[859], memory[858], memory[857], memory[856]},
        .ls2cmac_dat215       {memory[863], memory[862], memory[861], memory[860]},
        .ls2cmac_dat216       {memory[867], memory[866], memory[865], memory[864]},
        .ls2cmac_dat217       {memory[871], memory[870], memory[869], memory[868]},
        .ls2cmac_dat218       {memory[875], memory[874], memory[873], memory[872]},
        .ls2cmac_dat219       {memory[879], memory[878], memory[877], memory[876]},
        .ls2cmac_dat220       {memory[883], memory[882], memory[881], memory[880]},
        .ls2cmac_dat221       {memory[887], memory[886], memory[885], memory[884]},
        .ls2cmac_dat222       {memory[891], memory[890], memory[889], memory[888]},
        .ls2cmac_dat223       {memory[895], memory[894], memory[893], memory[892]},
        .ls2cmac_dat224       {memory[899], memory[898], memory[897], memory[896]},
        .ls2cmac_dat225       {memory[903], memory[902], memory[901], memory[900]},
        .ls2cmac_dat226       {memory[907], memory[906], memory[905], memory[904]},
        .ls2cmac_dat227       {memory[911], memory[910], memory[909], memory[908]},
        .ls2cmac_dat228       {memory[915], memory[914], memory[913], memory[912]},
        .ls2cmac_dat229       {memory[919], memory[918], memory[917], memory[916]},
        .ls2cmac_dat230       {memory[923], memory[922], memory[921], memory[920]},
        .ls2cmac_dat231       {memory[927], memory[926], memory[925], memory[924]},
        .ls2cmac_dat232       {memory[931], memory[930], memory[929], memory[928]},
        .ls2cmac_dat233       {memory[935], memory[934], memory[933], memory[932]},
        .ls2cmac_dat234       {memory[939], memory[938], memory[937], memory[936]},
        .ls2cmac_dat235       {memory[943], memory[942], memory[941], memory[940]},
        .ls2cmac_dat236       {memory[947], memory[946], memory[945], memory[944]},
        .ls2cmac_dat237       {memory[951], memory[950], memory[949], memory[948]},
        .ls2cmac_dat238       {memory[955], memory[954], memory[953], memory[952]},
        .ls2cmac_dat239       {memory[959], memory[958], memory[957], memory[956]},
        .ls2cmac_dat240       {memory[963], memory[962], memory[961], memory[960]},
        .ls2cmac_dat241       {memory[967], memory[966], memory[965], memory[964]},
        .ls2cmac_dat242       {memory[971], memory[970], memory[969], memory[968]},
        .ls2cmac_dat243       {memory[975], memory[974], memory[973], memory[972]},
        .ls2cmac_dat244       {memory[979], memory[978], memory[977], memory[976]},
        .ls2cmac_dat245       {memory[983], memory[982], memory[981], memory[980]},
        .ls2cmac_dat246       {memory[987], memory[986], memory[985], memory[984]},
        .ls2cmac_dat247       {memory[991], memory[990], memory[989], memory[988]},
        .ls2cmac_dat248       {memory[995], memory[994], memory[993], memory[992]},
        .ls2cmac_dat249       {memory[999], memory[998], memory[997], memory[996]},
        .ls2cmac_dat250       {memory[1003], memory[1002], memory[1001], memory[1000]},
        .ls2cmac_dat251       {memory[1007], memory[1006], memory[1005], memory[1004]},
        .ls2cmac_dat252       {memory[1011], memory[1010], memory[1009], memory[1008]},
        .ls2cmac_dat253       {memory[1015], memory[1014], memory[1013], memory[1012]},
        .ls2cmac_dat254       {memory[1019], memory[1018], memory[1017], memory[1016]},
        .ls2cmac_dat255       {memory[1023], memory[1022], memory[1021], memory[1020]},
        .ls2cmac_dat256       {memory[1027], memory[1026], memory[1025], memory[1024]},
        .ls2cmac_dat257       {memory[1031], memory[1030], memory[1029], memory[1028]},
        .ls2cmac_dat258       {memory[1035], memory[1034], memory[1033], memory[1032]},
        .ls2cmac_dat259       {memory[1039], memory[1038], memory[1037], memory[1036]},
        .ls2cmac_dat260       {memory[1043], memory[1042], memory[1041], memory[1040]},
        .ls2cmac_dat261       {memory[1047], memory[1046], memory[1045], memory[1044]},
        .ls2cmac_dat262       {memory[1051], memory[1050], memory[1049], memory[1048]},
        .ls2cmac_dat263       {memory[1055], memory[1054], memory[1053], memory[1052]},
        .ls2cmac_dat264       {memory[1059], memory[1058], memory[1057], memory[1056]},
        .ls2cmac_dat265       {memory[1063], memory[1062], memory[1061], memory[1060]},
        .ls2cmac_dat266       {memory[1067], memory[1066], memory[1065], memory[1064]},
        .ls2cmac_dat267       {memory[1071], memory[1070], memory[1069], memory[1068]},
        .ls2cmac_dat268       {memory[1075], memory[1074], memory[1073], memory[1072]},
        .ls2cmac_dat269       {memory[1079], memory[1078], memory[1077], memory[1076]},
        .ls2cmac_dat270       {memory[1083], memory[1082], memory[1081], memory[1080]},
        .ls2cmac_dat271       {memory[1087], memory[1086], memory[1085], memory[1084]},
        .ls2cmac_dat272       {memory[1091], memory[1090], memory[1089], memory[1088]},
        .ls2cmac_dat273       {memory[1095], memory[1094], memory[1093], memory[1092]},
        .ls2cmac_dat274       {memory[1099], memory[1098], memory[1097], memory[1096]},
        .ls2cmac_dat275       {memory[1103], memory[1102], memory[1101], memory[1100]},
        .ls2cmac_dat276       {memory[1107], memory[1106], memory[1105], memory[1104]},
        .ls2cmac_dat277       {memory[1111], memory[1110], memory[1109], memory[1108]},
        .ls2cmac_dat278       {memory[1115], memory[1114], memory[1113], memory[1112]},
        .ls2cmac_dat279       {memory[1119], memory[1118], memory[1117], memory[1116]},
        .ls2cmac_dat280       {memory[1123], memory[1122], memory[1121], memory[1120]},
        .ls2cmac_dat281       {memory[1127], memory[1126], memory[1125], memory[1124]},
        .ls2cmac_dat282       {memory[1131], memory[1130], memory[1129], memory[1128]},
        .ls2cmac_dat283       {memory[1135], memory[1134], memory[1133], memory[1132]},
        .ls2cmac_dat284       {memory[1139], memory[1138], memory[1137], memory[1136]},
        .ls2cmac_dat285       {memory[1143], memory[1142], memory[1141], memory[1140]},
        .ls2cmac_dat286       {memory[1147], memory[1146], memory[1145], memory[1144]},
        .ls2cmac_dat287       {memory[1151], memory[1150], memory[1149], memory[1148]},
        .ls2cmac_dat288       {memory[1155], memory[1154], memory[1153], memory[1152]},
        .ls2cmac_dat289       {memory[1159], memory[1158], memory[1157], memory[1156]},
        .ls2cmac_dat290       {memory[1163], memory[1162], memory[1161], memory[1160]},
        .ls2cmac_dat291       {memory[1167], memory[1166], memory[1165], memory[1164]},
        .ls2cmac_dat292       {memory[1171], memory[1170], memory[1169], memory[1168]},
        .ls2cmac_dat293       {memory[1175], memory[1174], memory[1173], memory[1172]},
        .ls2cmac_dat294       {memory[1179], memory[1178], memory[1177], memory[1176]},
        .ls2cmac_dat295       {memory[1183], memory[1182], memory[1181], memory[1180]},
        .ls2cmac_dat296       {memory[1187], memory[1186], memory[1185], memory[1184]},
        .ls2cmac_dat297       {memory[1191], memory[1190], memory[1189], memory[1188]},
        .ls2cmac_dat298       {memory[1195], memory[1194], memory[1193], memory[1192]},
        .ls2cmac_dat299       {memory[1199], memory[1198], memory[1197], memory[1196]},
        .ls2cmac_dat300       {memory[1203], memory[1202], memory[1201], memory[1200]},
        .ls2cmac_dat301       {memory[1207], memory[1206], memory[1205], memory[1204]},
        .ls2cmac_dat302       {memory[1211], memory[1210], memory[1209], memory[1208]},
        .ls2cmac_dat303       {memory[1215], memory[1214], memory[1213], memory[1212]},
        .ls2cmac_dat304       {memory[1219], memory[1218], memory[1217], memory[1216]},
        .ls2cmac_dat305       {memory[1223], memory[1222], memory[1221], memory[1220]},
        .ls2cmac_dat306       {memory[1227], memory[1226], memory[1225], memory[1224]},
        .ls2cmac_dat307       {memory[1231], memory[1230], memory[1229], memory[1228]},
        .ls2cmac_dat308       {memory[1235], memory[1234], memory[1233], memory[1232]},
        .ls2cmac_dat309       {memory[1239], memory[1238], memory[1237], memory[1236]},
        .ls2cmac_dat310       {memory[1243], memory[1242], memory[1241], memory[1240]},
        .ls2cmac_dat311       {memory[1247], memory[1246], memory[1245], memory[1244]},
        .ls2cmac_dat312       {memory[1251], memory[1250], memory[1249], memory[1248]},
        .ls2cmac_dat313       {memory[1255], memory[1254], memory[1253], memory[1252]},
        .ls2cmac_dat314       {memory[1259], memory[1258], memory[1257], memory[1256]},
        .ls2cmac_dat315       {memory[1263], memory[1262], memory[1261], memory[1260]},
        .ls2cmac_dat316       {memory[1267], memory[1266], memory[1265], memory[1264]},
        .ls2cmac_dat317       {memory[1271], memory[1270], memory[1269], memory[1268]},
        .ls2cmac_dat318       {memory[1275], memory[1274], memory[1273], memory[1272]},
        .ls2cmac_dat319       {memory[1279], memory[1278], memory[1277], memory[1276]},
        .ls2cmac_dat320       {memory[1283], memory[1282], memory[1281], memory[1280]},
        .ls2cmac_dat321       {memory[1287], memory[1286], memory[1285], memory[1284]},
        .ls2cmac_dat322       {memory[1291], memory[1290], memory[1289], memory[1288]},
        .ls2cmac_dat323       {memory[1295], memory[1294], memory[1293], memory[1292]},
        .ls2cmac_dat324       {memory[1299], memory[1298], memory[1297], memory[1296]},
        .ls2cmac_dat325       {memory[1303], memory[1302], memory[1301], memory[1300]},
        .ls2cmac_dat326       {memory[1307], memory[1306], memory[1305], memory[1304]},
        .ls2cmac_dat327       {memory[1311], memory[1310], memory[1309], memory[1308]},
        .ls2cmac_dat328       {memory[1315], memory[1314], memory[1313], memory[1312]},
        .ls2cmac_dat329       {memory[1319], memory[1318], memory[1317], memory[1316]},
        .ls2cmac_dat330       {memory[1323], memory[1322], memory[1321], memory[1320]},
        .ls2cmac_dat331       {memory[1327], memory[1326], memory[1325], memory[1324]},
        .ls2cmac_dat332       {memory[1331], memory[1330], memory[1329], memory[1328]},
        .ls2cmac_dat333       {memory[1335], memory[1334], memory[1333], memory[1332]},
        .ls2cmac_dat334       {memory[1339], memory[1338], memory[1337], memory[1336]},
        .ls2cmac_dat335       {memory[1343], memory[1342], memory[1341], memory[1340]},
        .ls2cmac_dat336       {memory[1347], memory[1346], memory[1345], memory[1344]},
        .ls2cmac_dat337       {memory[1351], memory[1350], memory[1349], memory[1348]},
        .ls2cmac_dat338       {memory[1355], memory[1354], memory[1353], memory[1352]},
        .ls2cmac_dat339       {memory[1359], memory[1358], memory[1357], memory[1356]},
        .ls2cmac_dat340       {memory[1363], memory[1362], memory[1361], memory[1360]},
        .ls2cmac_dat341       {memory[1367], memory[1366], memory[1365], memory[1364]},
        .ls2cmac_dat342       {memory[1371], memory[1370], memory[1369], memory[1368]},
        .ls2cmac_dat343       {memory[1375], memory[1374], memory[1373], memory[1372]},
        .ls2cmac_dat344       {memory[1379], memory[1378], memory[1377], memory[1376]},
        .ls2cmac_dat345       {memory[1383], memory[1382], memory[1381], memory[1380]},
        .ls2cmac_dat346       {memory[1387], memory[1386], memory[1385], memory[1384]},
        .ls2cmac_dat347       {memory[1391], memory[1390], memory[1389], memory[1388]},
        .ls2cmac_dat348       {memory[1395], memory[1394], memory[1393], memory[1392]},
        .ls2cmac_dat349       {memory[1399], memory[1398], memory[1397], memory[1396]},
        .ls2cmac_dat350       {memory[1403], memory[1402], memory[1401], memory[1400]},
        .ls2cmac_dat351       {memory[1407], memory[1406], memory[1405], memory[1404]},
        .ls2cmac_dat352       {memory[1411], memory[1410], memory[1409], memory[1408]},
        .ls2cmac_dat353       {memory[1415], memory[1414], memory[1413], memory[1412]},
        .ls2cmac_dat354       {memory[1419], memory[1418], memory[1417], memory[1416]},
        .ls2cmac_dat355       {memory[1423], memory[1422], memory[1421], memory[1420]},
        .ls2cmac_dat356       {memory[1427], memory[1426], memory[1425], memory[1424]},
        .ls2cmac_dat357       {memory[1431], memory[1430], memory[1429], memory[1428]},
        .ls2cmac_dat358       {memory[1435], memory[1434], memory[1433], memory[1432]},
        .ls2cmac_dat359       {memory[1439], memory[1438], memory[1437], memory[1436]},
        .ls2cmac_dat360       {memory[1443], memory[1442], memory[1441], memory[1440]},
        .ls2cmac_dat361       {memory[1447], memory[1446], memory[1445], memory[1444]},
        .ls2cmac_dat362       {memory[1451], memory[1450], memory[1449], memory[1448]},
        .ls2cmac_dat363       {memory[1455], memory[1454], memory[1453], memory[1452]},
        .ls2cmac_dat364       {memory[1459], memory[1458], memory[1457], memory[1456]},
        .ls2cmac_dat365       {memory[1463], memory[1462], memory[1461], memory[1460]},
        .ls2cmac_dat366       {memory[1467], memory[1466], memory[1465], memory[1464]},
        .ls2cmac_dat367       {memory[1471], memory[1470], memory[1469], memory[1468]},
        .ls2cmac_dat368       {memory[1475], memory[1474], memory[1473], memory[1472]},
        .ls2cmac_dat369       {memory[1479], memory[1478], memory[1477], memory[1476]},
        .ls2cmac_dat370       {memory[1483], memory[1482], memory[1481], memory[1480]},
        .ls2cmac_dat371       {memory[1487], memory[1486], memory[1485], memory[1484]},
        .ls2cmac_dat372       {memory[1491], memory[1490], memory[1489], memory[1488]},
        .ls2cmac_dat373       {memory[1495], memory[1494], memory[1493], memory[1492]},
        .ls2cmac_dat374       {memory[1499], memory[1498], memory[1497], memory[1496]},
        .ls2cmac_dat375       {memory[1503], memory[1502], memory[1501], memory[1500]},
        .ls2cmac_dat376       {memory[1507], memory[1506], memory[1505], memory[1504]},
        .ls2cmac_dat377       {memory[1511], memory[1510], memory[1509], memory[1508]},
        .ls2cmac_dat378       {memory[1515], memory[1514], memory[1513], memory[1512]},
        .ls2cmac_dat379       {memory[1519], memory[1518], memory[1517], memory[1516]},
        .ls2cmac_dat380       {memory[1523], memory[1522], memory[1521], memory[1520]},
        .ls2cmac_dat381       {memory[1527], memory[1526], memory[1525], memory[1524]},
        .ls2cmac_dat382       {memory[1531], memory[1530], memory[1529], memory[1528]},
        .ls2cmac_dat383       {memory[1535], memory[1534], memory[1533], memory[1532]},
        .ls2cmac_dat384       {memory[1539], memory[1538], memory[1537], memory[1536]},
        .ls2cmac_dat385       {memory[1543], memory[1542], memory[1541], memory[1540]},
        .ls2cmac_dat386       {memory[1547], memory[1546], memory[1545], memory[1544]},
        .ls2cmac_dat387       {memory[1551], memory[1550], memory[1549], memory[1548]},
        .ls2cmac_dat388       {memory[1555], memory[1554], memory[1553], memory[1552]},
        .ls2cmac_dat389       {memory[1559], memory[1558], memory[1557], memory[1556]},
        .ls2cmac_dat390       {memory[1563], memory[1562], memory[1561], memory[1560]},
        .ls2cmac_dat391       {memory[1567], memory[1566], memory[1565], memory[1564]},
        .ls2cmac_dat392       {memory[1571], memory[1570], memory[1569], memory[1568]},
        .ls2cmac_dat393       {memory[1575], memory[1574], memory[1573], memory[1572]},
        .ls2cmac_dat394       {memory[1579], memory[1578], memory[1577], memory[1576]},
        .ls2cmac_dat395       {memory[1583], memory[1582], memory[1581], memory[1580]},
        .ls2cmac_dat396       {memory[1587], memory[1586], memory[1585], memory[1584]},
        .ls2cmac_dat397       {memory[1591], memory[1590], memory[1589], memory[1588]},
        .ls2cmac_dat398       {memory[1595], memory[1594], memory[1593], memory[1592]},
        .ls2cmac_dat399       {memory[1599], memory[1598], memory[1597], memory[1596]},
        .ls2cmac_dat400       {memory[1603], memory[1602], memory[1601], memory[1600]},
        .ls2cmac_dat401       {memory[1607], memory[1606], memory[1605], memory[1604]},
        .ls2cmac_dat402       {memory[1611], memory[1610], memory[1609], memory[1608]},
        .ls2cmac_dat403       {memory[1615], memory[1614], memory[1613], memory[1612]},
        .ls2cmac_dat404       {memory[1619], memory[1618], memory[1617], memory[1616]},
        .ls2cmac_dat405       {memory[1623], memory[1622], memory[1621], memory[1620]},
        .ls2cmac_dat406       {memory[1627], memory[1626], memory[1625], memory[1624]},
        .ls2cmac_dat407       {memory[1631], memory[1630], memory[1629], memory[1628]},
        .ls2cmac_dat408       {memory[1635], memory[1634], memory[1633], memory[1632]},
        .ls2cmac_dat409       {memory[1639], memory[1638], memory[1637], memory[1636]},
        .ls2cmac_dat410       {memory[1643], memory[1642], memory[1641], memory[1640]},
        .ls2cmac_dat411       {memory[1647], memory[1646], memory[1645], memory[1644]},
        .ls2cmac_dat412       {memory[1651], memory[1650], memory[1649], memory[1648]},
        .ls2cmac_dat413       {memory[1655], memory[1654], memory[1653], memory[1652]},
        .ls2cmac_dat414       {memory[1659], memory[1658], memory[1657], memory[1656]},
        .ls2cmac_dat415       {memory[1663], memory[1662], memory[1661], memory[1660]},
        .ls2cmac_dat416       {memory[1667], memory[1666], memory[1665], memory[1664]},
        .ls2cmac_dat417       {memory[1671], memory[1670], memory[1669], memory[1668]},
        .ls2cmac_dat418       {memory[1675], memory[1674], memory[1673], memory[1672]},
        .ls2cmac_dat419       {memory[1679], memory[1678], memory[1677], memory[1676]},
        .ls2cmac_dat420       {memory[1683], memory[1682], memory[1681], memory[1680]},
        .ls2cmac_dat421       {memory[1687], memory[1686], memory[1685], memory[1684]},
        .ls2cmac_dat422       {memory[1691], memory[1690], memory[1689], memory[1688]},
        .ls2cmac_dat423       {memory[1695], memory[1694], memory[1693], memory[1692]},
        .ls2cmac_dat424       {memory[1699], memory[1698], memory[1697], memory[1696]},
        .ls2cmac_dat425       {memory[1703], memory[1702], memory[1701], memory[1700]},
        .ls2cmac_dat426       {memory[1707], memory[1706], memory[1705], memory[1704]},
        .ls2cmac_dat427       {memory[1711], memory[1710], memory[1709], memory[1708]},
        .ls2cmac_dat428       {memory[1715], memory[1714], memory[1713], memory[1712]},
        .ls2cmac_dat429       {memory[1719], memory[1718], memory[1717], memory[1716]},
        .ls2cmac_dat430       {memory[1723], memory[1722], memory[1721], memory[1720]},
        .ls2cmac_dat431       {memory[1727], memory[1726], memory[1725], memory[1724]},
        .ls2cmac_dat432       {memory[1731], memory[1730], memory[1729], memory[1728]},
        .ls2cmac_dat433       {memory[1735], memory[1734], memory[1733], memory[1732]},
        .ls2cmac_dat434       {memory[1739], memory[1738], memory[1737], memory[1736]},
        .ls2cmac_dat435       {memory[1743], memory[1742], memory[1741], memory[1740]},
        .ls2cmac_dat436       {memory[1747], memory[1746], memory[1745], memory[1744]},
        .ls2cmac_dat437       {memory[1751], memory[1750], memory[1749], memory[1748]},
        .ls2cmac_dat438       {memory[1755], memory[1754], memory[1753], memory[1752]},
        .ls2cmac_dat439       {memory[1759], memory[1758], memory[1757], memory[1756]},
        .ls2cmac_dat440       {memory[1763], memory[1762], memory[1761], memory[1760]},
        .ls2cmac_dat441       {memory[1767], memory[1766], memory[1765], memory[1764]},
        .ls2cmac_dat442       {memory[1771], memory[1770], memory[1769], memory[1768]},
        .ls2cmac_dat443       {memory[1775], memory[1774], memory[1773], memory[1772]},
        .ls2cmac_dat444       {memory[1779], memory[1778], memory[1777], memory[1776]},
        .ls2cmac_dat445       {memory[1783], memory[1782], memory[1781], memory[1780]},
        .ls2cmac_dat446       {memory[1787], memory[1786], memory[1785], memory[1784]},
        .ls2cmac_dat447       {memory[1791], memory[1790], memory[1789], memory[1788]},
        .ls2cmac_dat448       {memory[1795], memory[1794], memory[1793], memory[1792]},
        .ls2cmac_dat449       {memory[1799], memory[1798], memory[1797], memory[1796]},
        .ls2cmac_dat450       {memory[1803], memory[1802], memory[1801], memory[1800]},
        .ls2cmac_dat451       {memory[1807], memory[1806], memory[1805], memory[1804]},
        .ls2cmac_dat452       {memory[1811], memory[1810], memory[1809], memory[1808]},
        .ls2cmac_dat453       {memory[1815], memory[1814], memory[1813], memory[1812]},
        .ls2cmac_dat454       {memory[1819], memory[1818], memory[1817], memory[1816]},
        .ls2cmac_dat455       {memory[1823], memory[1822], memory[1821], memory[1820]},
        .ls2cmac_dat456       {memory[1827], memory[1826], memory[1825], memory[1824]},
        .ls2cmac_dat457       {memory[1831], memory[1830], memory[1829], memory[1828]},
        .ls2cmac_dat458       {memory[1835], memory[1834], memory[1833], memory[1832]},
        .ls2cmac_dat459       {memory[1839], memory[1838], memory[1837], memory[1836]},
        .ls2cmac_dat460       {memory[1843], memory[1842], memory[1841], memory[1840]},
        .ls2cmac_dat461       {memory[1847], memory[1846], memory[1845], memory[1844]},
        .ls2cmac_dat462       {memory[1851], memory[1850], memory[1849], memory[1848]},
        .ls2cmac_dat463       {memory[1855], memory[1854], memory[1853], memory[1852]},
        .ls2cmac_dat464       {memory[1859], memory[1858], memory[1857], memory[1856]},
        .ls2cmac_dat465       {memory[1863], memory[1862], memory[1861], memory[1860]},
        .ls2cmac_dat466       {memory[1867], memory[1866], memory[1865], memory[1864]},
        .ls2cmac_dat467       {memory[1871], memory[1870], memory[1869], memory[1868]},
        .ls2cmac_dat468       {memory[1875], memory[1874], memory[1873], memory[1872]},
        .ls2cmac_dat469       {memory[1879], memory[1878], memory[1877], memory[1876]},
        .ls2cmac_dat470       {memory[1883], memory[1882], memory[1881], memory[1880]},
        .ls2cmac_dat471       {memory[1887], memory[1886], memory[1885], memory[1884]},
        .ls2cmac_dat472       {memory[1891], memory[1890], memory[1889], memory[1888]},
        .ls2cmac_dat473       {memory[1895], memory[1894], memory[1893], memory[1892]},
        .ls2cmac_dat474       {memory[1899], memory[1898], memory[1897], memory[1896]},
        .ls2cmac_dat475       {memory[1903], memory[1902], memory[1901], memory[1900]},
        .ls2cmac_dat476       {memory[1907], memory[1906], memory[1905], memory[1904]},
        .ls2cmac_dat477       {memory[1911], memory[1910], memory[1909], memory[1908]},
        .ls2cmac_dat478       {memory[1915], memory[1914], memory[1913], memory[1912]},
        .ls2cmac_dat479       {memory[1919], memory[1918], memory[1917], memory[1916]},
        .ls2cmac_dat480       {memory[1923], memory[1922], memory[1921], memory[1920]},
        .ls2cmac_dat481       {memory[1927], memory[1926], memory[1925], memory[1924]},
        .ls2cmac_dat482       {memory[1931], memory[1930], memory[1929], memory[1928]},
        .ls2cmac_dat483       {memory[1935], memory[1934], memory[1933], memory[1932]},
        .ls2cmac_dat484       {memory[1939], memory[1938], memory[1937], memory[1936]},
        .ls2cmac_dat485       {memory[1943], memory[1942], memory[1941], memory[1940]},
        .ls2cmac_dat486       {memory[1947], memory[1946], memory[1945], memory[1944]},
        .ls2cmac_dat487       {memory[1951], memory[1950], memory[1949], memory[1948]},
        .ls2cmac_dat488       {memory[1955], memory[1954], memory[1953], memory[1952]},
        .ls2cmac_dat489       {memory[1959], memory[1958], memory[1957], memory[1956]},
        .ls2cmac_dat490       {memory[1963], memory[1962], memory[1961], memory[1960]},
        .ls2cmac_dat491       {memory[1967], memory[1966], memory[1965], memory[1964]},
        .ls2cmac_dat492       {memory[1971], memory[1970], memory[1969], memory[1968]},
        .ls2cmac_dat493       {memory[1975], memory[1974], memory[1973], memory[1972]},
        .ls2cmac_dat494       {memory[1979], memory[1978], memory[1977], memory[1976]},
        .ls2cmac_dat495       {memory[1983], memory[1982], memory[1981], memory[1980]},
        .ls2cmac_dat496       {memory[1987], memory[1986], memory[1985], memory[1984]},
        .ls2cmac_dat497       {memory[1991], memory[1990], memory[1989], memory[1988]},
        .ls2cmac_dat498       {memory[1995], memory[1994], memory[1993], memory[1992]},
        .ls2cmac_dat499       {memory[1999], memory[1998], memory[1997], memory[1996]},
        .ls2cmac_dat500       {memory[2003], memory[2002], memory[2001], memory[2000]},
        .ls2cmac_dat501       {memory[2007], memory[2006], memory[2005], memory[2004]},
        .ls2cmac_dat502       {memory[2011], memory[2010], memory[2009], memory[2008]},
        .ls2cmac_dat503       {memory[2015], memory[2014], memory[2013], memory[2012]},
        .ls2cmac_dat504       {memory[2019], memory[2018], memory[2017], memory[2016]},
        .ls2cmac_dat505       {memory[2023], memory[2022], memory[2021], memory[2020]},
        .ls2cmac_dat506       {memory[2027], memory[2026], memory[2025], memory[2024]},
        .ls2cmac_dat507       {memory[2031], memory[2030], memory[2029], memory[2028]},
        .ls2cmac_dat508       {memory[2035], memory[2034], memory[2033], memory[2032]},
        .ls2cmac_dat509       {memory[2039], memory[2038], memory[2037], memory[2036]},
        .ls2cmac_dat510       {memory[2043], memory[2042], memory[2041], memory[2040]},
        .ls2cmac_dat511       {memory[2047], memory[2046], memory[2045], memory[2044]},
        .ls2cmac_dat512       {memory[2051], memory[2050], memory[2049], memory[2048]},
        .ls2cmac_dat513       {memory[2055], memory[2054], memory[2053], memory[2052]},
        .ls2cmac_dat514       {memory[2059], memory[2058], memory[2057], memory[2056]},
        .ls2cmac_dat515       {memory[2063], memory[2062], memory[2061], memory[2060]},
        .ls2cmac_dat516       {memory[2067], memory[2066], memory[2065], memory[2064]},
        .ls2cmac_dat517       {memory[2071], memory[2070], memory[2069], memory[2068]},
        .ls2cmac_dat518       {memory[2075], memory[2074], memory[2073], memory[2072]},
        .ls2cmac_dat519       {memory[2079], memory[2078], memory[2077], memory[2076]},
        .ls2cmac_dat520       {memory[2083], memory[2082], memory[2081], memory[2080]},
        .ls2cmac_dat521       {memory[2087], memory[2086], memory[2085], memory[2084]},
        .ls2cmac_dat522       {memory[2091], memory[2090], memory[2089], memory[2088]},
        .ls2cmac_dat523       {memory[2095], memory[2094], memory[2093], memory[2092]},
        .ls2cmac_dat524       {memory[2099], memory[2098], memory[2097], memory[2096]},
        .ls2cmac_dat525       {memory[2103], memory[2102], memory[2101], memory[2100]},
        .ls2cmac_dat526       {memory[2107], memory[2106], memory[2105], memory[2104]},
        .ls2cmac_dat527       {memory[2111], memory[2110], memory[2109], memory[2108]},
        .ls2cmac_dat528       {memory[2115], memory[2114], memory[2113], memory[2112]},
        .ls2cmac_dat529       {memory[2119], memory[2118], memory[2117], memory[2116]},
        .ls2cmac_dat530       {memory[2123], memory[2122], memory[2121], memory[2120]},
        .ls2cmac_dat531       {memory[2127], memory[2126], memory[2125], memory[2124]},
        .ls2cmac_dat532       {memory[2131], memory[2130], memory[2129], memory[2128]},
        .ls2cmac_dat533       {memory[2135], memory[2134], memory[2133], memory[2132]},
        .ls2cmac_dat534       {memory[2139], memory[2138], memory[2137], memory[2136]},
        .ls2cmac_dat535       {memory[2143], memory[2142], memory[2141], memory[2140]},
        .ls2cmac_dat536       {memory[2147], memory[2146], memory[2145], memory[2144]},
        .ls2cmac_dat537       {memory[2151], memory[2150], memory[2149], memory[2148]},
        .ls2cmac_dat538       {memory[2155], memory[2154], memory[2153], memory[2152]},
        .ls2cmac_dat539       {memory[2159], memory[2158], memory[2157], memory[2156]},
        .ls2cmac_dat540       {memory[2163], memory[2162], memory[2161], memory[2160]},
        .ls2cmac_dat541       {memory[2167], memory[2166], memory[2165], memory[2164]},
        .ls2cmac_dat542       {memory[2171], memory[2170], memory[2169], memory[2168]},
        .ls2cmac_dat543       {memory[2175], memory[2174], memory[2173], memory[2172]},
        .ls2cmac_dat544       {memory[2179], memory[2178], memory[2177], memory[2176]},
        .ls2cmac_dat545       {memory[2183], memory[2182], memory[2181], memory[2180]},
        .ls2cmac_dat546       {memory[2187], memory[2186], memory[2185], memory[2184]},
        .ls2cmac_dat547       {memory[2191], memory[2190], memory[2189], memory[2188]},
        .ls2cmac_dat548       {memory[2195], memory[2194], memory[2193], memory[2192]},
        .ls2cmac_dat549       {memory[2199], memory[2198], memory[2197], memory[2196]},
        .ls2cmac_dat550       {memory[2203], memory[2202], memory[2201], memory[2200]},
        .ls2cmac_dat551       {memory[2207], memory[2206], memory[2205], memory[2204]},
        .ls2cmac_dat552       {memory[2211], memory[2210], memory[2209], memory[2208]},
        .ls2cmac_dat553       {memory[2215], memory[2214], memory[2213], memory[2212]},
        .ls2cmac_dat554       {memory[2219], memory[2218], memory[2217], memory[2216]},
        .ls2cmac_dat555       {memory[2223], memory[2222], memory[2221], memory[2220]},
        .ls2cmac_dat556       {memory[2227], memory[2226], memory[2225], memory[2224]},
        .ls2cmac_dat557       {memory[2231], memory[2230], memory[2229], memory[2228]},
        .ls2cmac_dat558       {memory[2235], memory[2234], memory[2233], memory[2232]},
        .ls2cmac_dat559       {memory[2239], memory[2238], memory[2237], memory[2236]},
        .ls2cmac_dat560       {memory[2243], memory[2242], memory[2241], memory[2240]},
        .ls2cmac_dat561       {memory[2247], memory[2246], memory[2245], memory[2244]},
        .ls2cmac_dat562       {memory[2251], memory[2250], memory[2249], memory[2248]},
        .ls2cmac_dat563       {memory[2255], memory[2254], memory[2253], memory[2252]},
        .ls2cmac_dat564       {memory[2259], memory[2258], memory[2257], memory[2256]},
        .ls2cmac_dat565       {memory[2263], memory[2262], memory[2261], memory[2260]},
        .ls2cmac_dat566       {memory[2267], memory[2266], memory[2265], memory[2264]},
        .ls2cmac_dat567       {memory[2271], memory[2270], memory[2269], memory[2268]},
        .ls2cmac_dat568       {memory[2275], memory[2274], memory[2273], memory[2272]},
        .ls2cmac_dat569       {memory[2279], memory[2278], memory[2277], memory[2276]},
        .ls2cmac_dat570       {memory[2283], memory[2282], memory[2281], memory[2280]},
        .ls2cmac_dat571       {memory[2287], memory[2286], memory[2285], memory[2284]},
        .ls2cmac_dat572       {memory[2291], memory[2290], memory[2289], memory[2288]},
        .ls2cmac_dat573       {memory[2295], memory[2294], memory[2293], memory[2292]},
        .ls2cmac_dat574       {memory[2299], memory[2298], memory[2297], memory[2296]},
        .ls2cmac_dat575       {memory[2303], memory[2302], memory[2301], memory[2300]},
        .ls2cmac_dat576       {memory[2307], memory[2306], memory[2305], memory[2304]},
        .ls2cmac_dat577       {memory[2311], memory[2310], memory[2309], memory[2308]},
        .ls2cmac_dat578       {memory[2315], memory[2314], memory[2313], memory[2312]},
        .ls2cmac_dat579       {memory[2319], memory[2318], memory[2317], memory[2316]},
        .ls2cmac_dat580       {memory[2323], memory[2322], memory[2321], memory[2320]},
        .ls2cmac_dat581       {memory[2327], memory[2326], memory[2325], memory[2324]},
        .ls2cmac_dat582       {memory[2331], memory[2330], memory[2329], memory[2328]},
        .ls2cmac_dat583       {memory[2335], memory[2334], memory[2333], memory[2332]},
        .ls2cmac_dat584       {memory[2339], memory[2338], memory[2337], memory[2336]},
        .ls2cmac_dat585       {memory[2343], memory[2342], memory[2341], memory[2340]},
        .ls2cmac_dat586       {memory[2347], memory[2346], memory[2345], memory[2344]},
        .ls2cmac_dat587       {memory[2351], memory[2350], memory[2349], memory[2348]},
        .ls2cmac_dat588       {memory[2355], memory[2354], memory[2353], memory[2352]},
        .ls2cmac_dat589       {memory[2359], memory[2358], memory[2357], memory[2356]},
        .ls2cmac_dat590       {memory[2363], memory[2362], memory[2361], memory[2360]},
        .ls2cmac_dat591       {memory[2367], memory[2366], memory[2365], memory[2364]},
        .ls2cmac_dat592       {memory[2371], memory[2370], memory[2369], memory[2368]},
        .ls2cmac_dat593       {memory[2375], memory[2374], memory[2373], memory[2372]},
        .ls2cmac_dat594       {memory[2379], memory[2378], memory[2377], memory[2376]},
        .ls2cmac_dat595       {memory[2383], memory[2382], memory[2381], memory[2380]},
        .ls2cmac_dat596       {memory[2387], memory[2386], memory[2385], memory[2384]},
        .ls2cmac_dat597       {memory[2391], memory[2390], memory[2389], memory[2388]},
        .ls2cmac_dat598       {memory[2395], memory[2394], memory[2393], memory[2392]},
        .ls2cmac_dat599       {memory[2399], memory[2398], memory[2397], memory[2396]},
        .ls2cmac_dat600       {memory[2403], memory[2402], memory[2401], memory[2400]},
        .ls2cmac_dat601       {memory[2407], memory[2406], memory[2405], memory[2404]},
        .ls2cmac_dat602       {memory[2411], memory[2410], memory[2409], memory[2408]},
        .ls2cmac_dat603       {memory[2415], memory[2414], memory[2413], memory[2412]},
        .ls2cmac_dat604       {memory[2419], memory[2418], memory[2417], memory[2416]},
        .ls2cmac_dat605       {memory[2423], memory[2422], memory[2421], memory[2420]},
        .ls2cmac_dat606       {memory[2427], memory[2426], memory[2425], memory[2424]},
        .ls2cmac_dat607       {memory[2431], memory[2430], memory[2429], memory[2428]},
        .ls2cmac_dat608       {memory[2435], memory[2434], memory[2433], memory[2432]},
        .ls2cmac_dat609       {memory[2439], memory[2438], memory[2437], memory[2436]},
        .ls2cmac_dat610       {memory[2443], memory[2442], memory[2441], memory[2440]},
        .ls2cmac_dat611       {memory[2447], memory[2446], memory[2445], memory[2444]},
        .ls2cmac_dat612       {memory[2451], memory[2450], memory[2449], memory[2448]},
        .ls2cmac_dat613       {memory[2455], memory[2454], memory[2453], memory[2452]},
        .ls2cmac_dat614       {memory[2459], memory[2458], memory[2457], memory[2456]},
        .ls2cmac_dat615       {memory[2463], memory[2462], memory[2461], memory[2460]},
        .ls2cmac_dat616       {memory[2467], memory[2466], memory[2465], memory[2464]},
        .ls2cmac_dat617       {memory[2471], memory[2470], memory[2469], memory[2468]},
        .ls2cmac_dat618       {memory[2475], memory[2474], memory[2473], memory[2472]},
        .ls2cmac_dat619       {memory[2479], memory[2478], memory[2477], memory[2476]},
        .ls2cmac_dat620       {memory[2483], memory[2482], memory[2481], memory[2480]},
        .ls2cmac_dat621       {memory[2487], memory[2486], memory[2485], memory[2484]},
        .ls2cmac_dat622       {memory[2491], memory[2490], memory[2489], memory[2488]},
        .ls2cmac_dat623       {memory[2495], memory[2494], memory[2493], memory[2492]},
        .ls2cmac_dat624       {memory[2499], memory[2498], memory[2497], memory[2496]},
        .ls2cmac_dat625       {memory[2503], memory[2502], memory[2501], memory[2500]},
        .ls2cmac_dat626       {memory[2507], memory[2506], memory[2505], memory[2504]},
        .ls2cmac_dat627       {memory[2511], memory[2510], memory[2509], memory[2508]},
        .ls2cmac_dat628       {memory[2515], memory[2514], memory[2513], memory[2512]},
        .ls2cmac_dat629       {memory[2519], memory[2518], memory[2517], memory[2516]},
        .ls2cmac_dat630       {memory[2523], memory[2522], memory[2521], memory[2520]},
        .ls2cmac_dat631       {memory[2527], memory[2526], memory[2525], memory[2524]},
        .ls2cmac_dat632       {memory[2531], memory[2530], memory[2529], memory[2528]},
        .ls2cmac_dat633       {memory[2535], memory[2534], memory[2533], memory[2532]},
        .ls2cmac_dat634       {memory[2539], memory[2538], memory[2537], memory[2536]},
        .ls2cmac_dat635       {memory[2543], memory[2542], memory[2541], memory[2540]},
        .ls2cmac_dat636       {memory[2547], memory[2546], memory[2545], memory[2544]},
        .ls2cmac_dat637       {memory[2551], memory[2550], memory[2549], memory[2548]},
        .ls2cmac_dat638       {memory[2555], memory[2554], memory[2553], memory[2552]},
        .ls2cmac_dat639       {memory[2559], memory[2558], memory[2557], memory[2556]},
        .ls2cmac_dat640       {memory[2563], memory[2562], memory[2561], memory[2560]},
        .ls2cmac_dat641       {memory[2567], memory[2566], memory[2565], memory[2564]},
        .ls2cmac_dat642       {memory[2571], memory[2570], memory[2569], memory[2568]},
        .ls2cmac_dat643       {memory[2575], memory[2574], memory[2573], memory[2572]},
        .ls2cmac_dat644       {memory[2579], memory[2578], memory[2577], memory[2576]},
        .ls2cmac_dat645       {memory[2583], memory[2582], memory[2581], memory[2580]},
        .ls2cmac_dat646       {memory[2587], memory[2586], memory[2585], memory[2584]},
        .ls2cmac_dat647       {memory[2591], memory[2590], memory[2589], memory[2588]},
        .ls2cmac_dat648       {memory[2595], memory[2594], memory[2593], memory[2592]},
        .ls2cmac_dat649       {memory[2599], memory[2598], memory[2597], memory[2596]},
        .ls2cmac_dat650       {memory[2603], memory[2602], memory[2601], memory[2600]},
        .ls2cmac_dat651       {memory[2607], memory[2606], memory[2605], memory[2604]},
        .ls2cmac_dat652       {memory[2611], memory[2610], memory[2609], memory[2608]},
        .ls2cmac_dat653       {memory[2615], memory[2614], memory[2613], memory[2612]},
        .ls2cmac_dat654       {memory[2619], memory[2618], memory[2617], memory[2616]},
        .ls2cmac_dat655       {memory[2623], memory[2622], memory[2621], memory[2620]},
        .ls2cmac_dat656       {memory[2627], memory[2626], memory[2625], memory[2624]},
        .ls2cmac_dat657       {memory[2631], memory[2630], memory[2629], memory[2628]},
        .ls2cmac_dat658       {memory[2635], memory[2634], memory[2633], memory[2632]},
        .ls2cmac_dat659       {memory[2639], memory[2638], memory[2637], memory[2636]},
        .ls2cmac_dat660       {memory[2643], memory[2642], memory[2641], memory[2640]},
        .ls2cmac_dat661       {memory[2647], memory[2646], memory[2645], memory[2644]},
        .ls2cmac_dat662       {memory[2651], memory[2650], memory[2649], memory[2648]},
        .ls2cmac_dat663       {memory[2655], memory[2654], memory[2653], memory[2652]},
        .ls2cmac_dat664       {memory[2659], memory[2658], memory[2657], memory[2656]},
        .ls2cmac_dat665       {memory[2663], memory[2662], memory[2661], memory[2660]},
        .ls2cmac_dat666       {memory[2667], memory[2666], memory[2665], memory[2664]},
        .ls2cmac_dat667       {memory[2671], memory[2670], memory[2669], memory[2668]},
        .ls2cmac_dat668       {memory[2675], memory[2674], memory[2673], memory[2672]},
        .ls2cmac_dat669       {memory[2679], memory[2678], memory[2677], memory[2676]},
        .ls2cmac_dat670       {memory[2683], memory[2682], memory[2681], memory[2680]},
        .ls2cmac_dat671       {memory[2687], memory[2686], memory[2685], memory[2684]},
        .ls2cmac_dat672       {memory[2691], memory[2690], memory[2689], memory[2688]},
        .ls2cmac_dat673       {memory[2695], memory[2694], memory[2693], memory[2692]},
        .ls2cmac_dat674       {memory[2699], memory[2698], memory[2697], memory[2696]},
        .ls2cmac_dat675       {memory[2703], memory[2702], memory[2701], memory[2700]},
        .ls2cmac_dat676       {memory[2707], memory[2706], memory[2705], memory[2704]},
        .ls2cmac_dat677       {memory[2711], memory[2710], memory[2709], memory[2708]},
        .ls2cmac_dat678       {memory[2715], memory[2714], memory[2713], memory[2712]},
        .ls2cmac_dat679       {memory[2719], memory[2718], memory[2717], memory[2716]},
        .ls2cmac_dat680       {memory[2723], memory[2722], memory[2721], memory[2720]},
        .ls2cmac_dat681       {memory[2727], memory[2726], memory[2725], memory[2724]},
        .ls2cmac_dat682       {memory[2731], memory[2730], memory[2729], memory[2728]},
        .ls2cmac_dat683       {memory[2735], memory[2734], memory[2733], memory[2732]},
        .ls2cmac_dat684       {memory[2739], memory[2738], memory[2737], memory[2736]},
        .ls2cmac_dat685       {memory[2743], memory[2742], memory[2741], memory[2740]},
        .ls2cmac_dat686       {memory[2747], memory[2746], memory[2745], memory[2744]},
        .ls2cmac_dat687       {memory[2751], memory[2750], memory[2749], memory[2748]},
        .ls2cmac_dat688       {memory[2755], memory[2754], memory[2753], memory[2752]},
        .ls2cmac_dat689       {memory[2759], memory[2758], memory[2757], memory[2756]},
        .ls2cmac_dat690       {memory[2763], memory[2762], memory[2761], memory[2760]},
        .ls2cmac_dat691       {memory[2767], memory[2766], memory[2765], memory[2764]},
        .ls2cmac_dat692       {memory[2771], memory[2770], memory[2769], memory[2768]},
        .ls2cmac_dat693       {memory[2775], memory[2774], memory[2773], memory[2772]},
        .ls2cmac_dat694       {memory[2779], memory[2778], memory[2777], memory[2776]},
        .ls2cmac_dat695       {memory[2783], memory[2782], memory[2781], memory[2780]},
        .ls2cmac_dat696       {memory[2787], memory[2786], memory[2785], memory[2784]},
        .ls2cmac_dat697       {memory[2791], memory[2790], memory[2789], memory[2788]},
        .ls2cmac_dat698       {memory[2795], memory[2794], memory[2793], memory[2792]},
        .ls2cmac_dat699       {memory[2799], memory[2798], memory[2797], memory[2796]},
        .ls2cmac_dat700       {memory[2803], memory[2802], memory[2801], memory[2800]},
        .ls2cmac_dat701       {memory[2807], memory[2806], memory[2805], memory[2804]},
        .ls2cmac_dat702       {memory[2811], memory[2810], memory[2809], memory[2808]},
        .ls2cmac_dat703       {memory[2815], memory[2814], memory[2813], memory[2812]},
        .ls2cmac_dat704       {memory[2819], memory[2818], memory[2817], memory[2816]},
        .ls2cmac_dat705       {memory[2823], memory[2822], memory[2821], memory[2820]},
        .ls2cmac_dat706       {memory[2827], memory[2826], memory[2825], memory[2824]},
        .ls2cmac_dat707       {memory[2831], memory[2830], memory[2829], memory[2828]},
        .ls2cmac_dat708       {memory[2835], memory[2834], memory[2833], memory[2832]},
        .ls2cmac_dat709       {memory[2839], memory[2838], memory[2837], memory[2836]},
        .ls2cmac_dat710       {memory[2843], memory[2842], memory[2841], memory[2840]},
        .ls2cmac_dat711       {memory[2847], memory[2846], memory[2845], memory[2844]},
        .ls2cmac_dat712       {memory[2851], memory[2850], memory[2849], memory[2848]},
        .ls2cmac_dat713       {memory[2855], memory[2854], memory[2853], memory[2852]},
        .ls2cmac_dat714       {memory[2859], memory[2858], memory[2857], memory[2856]},
        .ls2cmac_dat715       {memory[2863], memory[2862], memory[2861], memory[2860]},
        .ls2cmac_dat716       {memory[2867], memory[2866], memory[2865], memory[2864]},
        .ls2cmac_dat717       {memory[2871], memory[2870], memory[2869], memory[2868]},
        .ls2cmac_dat718       {memory[2875], memory[2874], memory[2873], memory[2872]},
        .ls2cmac_dat719       {memory[2879], memory[2878], memory[2877], memory[2876]},
        .ls2cmac_dat720       {memory[2883], memory[2882], memory[2881], memory[2880]},
        .ls2cmac_dat721       {memory[2887], memory[2886], memory[2885], memory[2884]},
        .ls2cmac_dat722       {memory[2891], memory[2890], memory[2889], memory[2888]},
        .ls2cmac_dat723       {memory[2895], memory[2894], memory[2893], memory[2892]},
        .ls2cmac_dat724       {memory[2899], memory[2898], memory[2897], memory[2896]},
        .ls2cmac_dat725       {memory[2903], memory[2902], memory[2901], memory[2900]},
        .ls2cmac_dat726       {memory[2907], memory[2906], memory[2905], memory[2904]},
        .ls2cmac_dat727       {memory[2911], memory[2910], memory[2909], memory[2908]},
        .ls2cmac_dat728       {memory[2915], memory[2914], memory[2913], memory[2912]},
        .ls2cmac_dat729       {memory[2919], memory[2918], memory[2917], memory[2916]},
        .ls2cmac_dat730       {memory[2923], memory[2922], memory[2921], memory[2920]},
        .ls2cmac_dat731       {memory[2927], memory[2926], memory[2925], memory[2924]},
        .ls2cmac_dat732       {memory[2931], memory[2930], memory[2929], memory[2928]},
        .ls2cmac_dat733       {memory[2935], memory[2934], memory[2933], memory[2932]},
        .ls2cmac_dat734       {memory[2939], memory[2938], memory[2937], memory[2936]},
        .ls2cmac_dat735       {memory[2943], memory[2942], memory[2941], memory[2940]},
        .ls2cmac_dat736       {memory[2947], memory[2946], memory[2945], memory[2944]},
        .ls2cmac_dat737       {memory[2951], memory[2950], memory[2949], memory[2948]},
        .ls2cmac_dat738       {memory[2955], memory[2954], memory[2953], memory[2952]},
        .ls2cmac_dat739       {memory[2959], memory[2958], memory[2957], memory[2956]},
        .ls2cmac_dat740       {memory[2963], memory[2962], memory[2961], memory[2960]},
        .ls2cmac_dat741       {memory[2967], memory[2966], memory[2965], memory[2964]},
        .ls2cmac_dat742       {memory[2971], memory[2970], memory[2969], memory[2968]},
        .ls2cmac_dat743       {memory[2975], memory[2974], memory[2973], memory[2972]},
        .ls2cmac_dat744       {memory[2979], memory[2978], memory[2977], memory[2976]},
        .ls2cmac_dat745       {memory[2983], memory[2982], memory[2981], memory[2980]},
        .ls2cmac_dat746       {memory[2987], memory[2986], memory[2985], memory[2984]},
        .ls2cmac_dat747       {memory[2991], memory[2990], memory[2989], memory[2988]},
        .ls2cmac_dat748       {memory[2995], memory[2994], memory[2993], memory[2992]},
        .ls2cmac_dat749       {memory[2999], memory[2998], memory[2997], memory[2996]},
        .ls2cmac_dat750       {memory[3003], memory[3002], memory[3001], memory[3000]},
        .ls2cmac_dat751       {memory[3007], memory[3006], memory[3005], memory[3004]},
        .ls2cmac_dat752       {memory[3011], memory[3010], memory[3009], memory[3008]},
        .ls2cmac_dat753       {memory[3015], memory[3014], memory[3013], memory[3012]},
        .ls2cmac_dat754       {memory[3019], memory[3018], memory[3017], memory[3016]},
        .ls2cmac_dat755       {memory[3023], memory[3022], memory[3021], memory[3020]},
        .ls2cmac_dat756       {memory[3027], memory[3026], memory[3025], memory[3024]},
        .ls2cmac_dat757       {memory[3031], memory[3030], memory[3029], memory[3028]},
        .ls2cmac_dat758       {memory[3035], memory[3034], memory[3033], memory[3032]},
        .ls2cmac_dat759       {memory[3039], memory[3038], memory[3037], memory[3036]},
        .ls2cmac_dat760       {memory[3043], memory[3042], memory[3041], memory[3040]},
        .ls2cmac_dat761       {memory[3047], memory[3046], memory[3045], memory[3044]},
        .ls2cmac_dat762       {memory[3051], memory[3050], memory[3049], memory[3048]},
        .ls2cmac_dat763       {memory[3055], memory[3054], memory[3053], memory[3052]},
        .ls2cmac_dat764       {memory[3059], memory[3058], memory[3057], memory[3056]},
        .ls2cmac_dat765       {memory[3063], memory[3062], memory[3061], memory[3060]},
        .ls2cmac_dat766       {memory[3067], memory[3066], memory[3065], memory[3064]},
        .ls2cmac_dat767       {memory[3071], memory[3070], memory[3069], memory[3068]},
        .ls2cmac_dat768       {memory[3075], memory[3074], memory[3073], memory[3072]},
        .ls2cmac_dat769       {memory[3079], memory[3078], memory[3077], memory[3076]},
        .ls2cmac_dat770       {memory[3083], memory[3082], memory[3081], memory[3080]},
        .ls2cmac_dat771       {memory[3087], memory[3086], memory[3085], memory[3084]},
        .ls2cmac_dat772       {memory[3091], memory[3090], memory[3089], memory[3088]},
        .ls2cmac_dat773       {memory[3095], memory[3094], memory[3093], memory[3092]},
        .ls2cmac_dat774       {memory[3099], memory[3098], memory[3097], memory[3096]},
        .ls2cmac_dat775       {memory[3103], memory[3102], memory[3101], memory[3100]},
        .ls2cmac_dat776       {memory[3107], memory[3106], memory[3105], memory[3104]},
        .ls2cmac_dat777       {memory[3111], memory[3110], memory[3109], memory[3108]},
        .ls2cmac_dat778       {memory[3115], memory[3114], memory[3113], memory[3112]},
        .ls2cmac_dat779       {memory[3119], memory[3118], memory[3117], memory[3116]},
        .ls2cmac_dat780       {memory[3123], memory[3122], memory[3121], memory[3120]},
        .ls2cmac_dat781       {memory[3127], memory[3126], memory[3125], memory[3124]},
        .ls2cmac_dat782       {memory[3131], memory[3130], memory[3129], memory[3128]},
        .ls2cmac_dat783       {memory[3135], memory[3134], memory[3133], memory[3132]},
        .ls2cmac_dat_size     data_size,
        .ls2cmac_wt0       {memory[3139], memory[3138], memory[3137], memory[3136]},
        .ls2cmac_wt1       {memory[3143], memory[3142], memory[3141], memory[3140]},
        .ls2cmac_wt2       {memory[3147], memory[3146], memory[3145], memory[3144]},
        .ls2cmac_wt3       {memory[3151], memory[3150], memory[3149], memory[3148]},
        .ls2cmac_wt4       {memory[3155], memory[3154], memory[3153], memory[3152]},
        .ls2cmac_wt5       {memory[3159], memory[3158], memory[3157], memory[3156]},
        .ls2cmac_wt6       {memory[3163], memory[3162], memory[3161], memory[3160]},
        .ls2cmac_wt7       {memory[3167], memory[3166], memory[3165], memory[3164]},
        .ls2cmac_wt8       {memory[3171], memory[3170], memory[3169], memory[3168]},
        .ls2cmac_wt9       {memory[3175], memory[3174], memory[3173], memory[3172]},
        .ls2cmac_wt10       {memory[3179], memory[3178], memory[3177], memory[3176]},
        .ls2cmac_wt11       {memory[3183], memory[3182], memory[3181], memory[3180]},
        .ls2cmac_wt12       {memory[3187], memory[3186], memory[3185], memory[3184]},
        .ls2cmac_wt13       {memory[3191], memory[3190], memory[3189], memory[3188]},
        .ls2cmac_wt14       {memory[3195], memory[3194], memory[3193], memory[3192]},
        .ls2cmac_wt15       {memory[3199], memory[3198], memory[3197], memory[3196]},
        .ls2cmac_wt16       {memory[3203], memory[3202], memory[3201], memory[3200]},
        .ls2cmac_wt17       {memory[3207], memory[3206], memory[3205], memory[3204]},
        .ls2cmac_wt18       {memory[3211], memory[3210], memory[3209], memory[3208]},
        .ls2cmac_wt19       {memory[3215], memory[3214], memory[3213], memory[3212]},
        .ls2cmac_wt20       {memory[3219], memory[3218], memory[3217], memory[3216]},
        .ls2cmac_wt21       {memory[3223], memory[3222], memory[3221], memory[3220]},
        .ls2cmac_wt22       {memory[3227], memory[3226], memory[3225], memory[3224]},
        .ls2cmac_wt23       {memory[3231], memory[3230], memory[3229], memory[3228]},
        .ls2cmac_wt24       {memory[3235], memory[3234], memory[3233], memory[3232]},
        .ls2cmac_wt_size        weight_size);


endmodule
