// ytydla_conv.sv

`include "ytydla_define.svh"


module ytydla_conv2d(ytydla_core_clk,
                     ytydla_core_rst_n,
                        ls2cmac_dat0,
                        ls2cmac_dat1,
                        ls2cmac_dat2,
                        ls2cmac_dat3,
                        ls2cmac_dat4,
                        ls2cmac_dat5,
                        ls2cmac_dat6,
                        ls2cmac_dat7,
                        ls2cmac_dat8,
                        ls2cmac_dat9,
                        ls2cmac_dat10,
                        ls2cmac_dat11,
                        ls2cmac_dat12,
                        ls2cmac_dat13,
                        ls2cmac_dat14,
                        ls2cmac_dat15,
                        ls2cmac_dat16,
                        ls2cmac_dat17,
                        ls2cmac_dat18,
                        ls2cmac_dat19,
                        ls2cmac_dat20,
                        ls2cmac_dat21,
                        ls2cmac_dat22,
                        ls2cmac_dat23,
                        ls2cmac_dat24,
                        ls2cmac_dat25,
                        ls2cmac_dat26,
                        ls2cmac_dat27,
                        ls2cmac_dat28,
                        ls2cmac_dat29,
                        ls2cmac_dat30,
                        ls2cmac_dat31,
                        ls2cmac_dat32,
                        ls2cmac_dat33,
                        ls2cmac_dat34,
                        ls2cmac_dat35,
                        ls2cmac_dat36,
                        ls2cmac_dat37,
                        ls2cmac_dat38,
                        ls2cmac_dat39,
                        ls2cmac_dat40,
                        ls2cmac_dat41,
                        ls2cmac_dat42,
                        ls2cmac_dat43,
                        ls2cmac_dat44,
                        ls2cmac_dat45,
                        ls2cmac_dat46,
                        ls2cmac_dat47,
                        ls2cmac_dat48,
                        ls2cmac_dat49,
                        ls2cmac_dat50,
                        ls2cmac_dat51,
                        ls2cmac_dat52,
                        ls2cmac_dat53,
                        ls2cmac_dat54,
                        ls2cmac_dat55,
                        ls2cmac_dat56,
                        ls2cmac_dat57,
                        ls2cmac_dat58,
                        ls2cmac_dat59,
                        ls2cmac_dat60,
                        ls2cmac_dat61,
                        ls2cmac_dat62,
                        ls2cmac_dat63,
                        ls2cmac_dat64,
                        ls2cmac_dat65,
                        ls2cmac_dat66,
                        ls2cmac_dat67,
                        ls2cmac_dat68,
                        ls2cmac_dat69,
                        ls2cmac_dat70,
                        ls2cmac_dat71,
                        ls2cmac_dat72,
                        ls2cmac_dat73,
                        ls2cmac_dat74,
                        ls2cmac_dat75,
                        ls2cmac_dat76,
                        ls2cmac_dat77,
                        ls2cmac_dat78,
                        ls2cmac_dat79,
                        ls2cmac_dat80,
                        ls2cmac_dat81,
                        ls2cmac_dat82,
                        ls2cmac_dat83,
                        ls2cmac_dat84,
                        ls2cmac_dat85,
                        ls2cmac_dat86,
                        ls2cmac_dat87,
                        ls2cmac_dat88,
                        ls2cmac_dat89,
                        ls2cmac_dat90,
                        ls2cmac_dat91,
                        ls2cmac_dat92,
                        ls2cmac_dat93,
                        ls2cmac_dat94,
                        ls2cmac_dat95,
                        ls2cmac_dat96,
                        ls2cmac_dat97,
                        ls2cmac_dat98,
                        ls2cmac_dat99,
                        ls2cmac_dat100,
                        ls2cmac_dat101,
                        ls2cmac_dat102,
                        ls2cmac_dat103,
                        ls2cmac_dat104,
                        ls2cmac_dat105,
                        ls2cmac_dat106,
                        ls2cmac_dat107,
                        ls2cmac_dat108,
                        ls2cmac_dat109,
                        ls2cmac_dat110,
                        ls2cmac_dat111,
                        ls2cmac_dat112,
                        ls2cmac_dat113,
                        ls2cmac_dat114,
                        ls2cmac_dat115,
                        ls2cmac_dat116,
                        ls2cmac_dat117,
                        ls2cmac_dat118,
                        ls2cmac_dat119,
                        ls2cmac_dat120,
                        ls2cmac_dat121,
                        ls2cmac_dat122,
                        ls2cmac_dat123,
                        ls2cmac_dat124,
                        ls2cmac_dat125,
                        ls2cmac_dat126,
                        ls2cmac_dat127,
                        ls2cmac_dat128,
                        ls2cmac_dat129,
                        ls2cmac_dat130,
                        ls2cmac_dat131,
                        ls2cmac_dat132,
                        ls2cmac_dat133,
                        ls2cmac_dat134,
                        ls2cmac_dat135,
                        ls2cmac_dat136,
                        ls2cmac_dat137,
                        ls2cmac_dat138,
                        ls2cmac_dat139,
                        ls2cmac_dat140,
                        ls2cmac_dat141,
                        ls2cmac_dat142,
                        ls2cmac_dat143,
                        ls2cmac_dat144,
                        ls2cmac_dat145,
                        ls2cmac_dat146,
                        ls2cmac_dat147,
                        ls2cmac_dat148,
                        ls2cmac_dat149,
                        ls2cmac_dat150,
                        ls2cmac_dat151,
                        ls2cmac_dat152,
                        ls2cmac_dat153,
                        ls2cmac_dat154,
                        ls2cmac_dat155,
                        ls2cmac_dat156,
                        ls2cmac_dat157,
                        ls2cmac_dat158,
                        ls2cmac_dat159,
                        ls2cmac_dat160,
                        ls2cmac_dat161,
                        ls2cmac_dat162,
                        ls2cmac_dat163,
                        ls2cmac_dat164,
                        ls2cmac_dat165,
                        ls2cmac_dat166,
                        ls2cmac_dat167,
                        ls2cmac_dat168,
                        ls2cmac_dat169,
                        ls2cmac_dat170,
                        ls2cmac_dat171,
                        ls2cmac_dat172,
                        ls2cmac_dat173,
                        ls2cmac_dat174,
                        ls2cmac_dat175,
                        ls2cmac_dat176,
                        ls2cmac_dat177,
                        ls2cmac_dat178,
                        ls2cmac_dat179,
                        ls2cmac_dat180,
                        ls2cmac_dat181,
                        ls2cmac_dat182,
                        ls2cmac_dat183,
                        ls2cmac_dat184,
                        ls2cmac_dat185,
                        ls2cmac_dat186,
                        ls2cmac_dat187,
                        ls2cmac_dat188,
                        ls2cmac_dat189,
                        ls2cmac_dat190,
                        ls2cmac_dat191,
                        ls2cmac_dat192,
                        ls2cmac_dat193,
                        ls2cmac_dat194,
                        ls2cmac_dat195,
                        ls2cmac_dat196,
                        ls2cmac_dat197,
                        ls2cmac_dat198,
                        ls2cmac_dat199,
                        ls2cmac_dat200,
                        ls2cmac_dat201,
                        ls2cmac_dat202,
                        ls2cmac_dat203,
                        ls2cmac_dat204,
                        ls2cmac_dat205,
                        ls2cmac_dat206,
                        ls2cmac_dat207,
                        ls2cmac_dat208,
                        ls2cmac_dat209,
                        ls2cmac_dat210,
                        ls2cmac_dat211,
                        ls2cmac_dat212,
                        ls2cmac_dat213,
                        ls2cmac_dat214,
                        ls2cmac_dat215,
                        ls2cmac_dat216,
                        ls2cmac_dat217,
                        ls2cmac_dat218,
                        ls2cmac_dat219,
                        ls2cmac_dat220,
                        ls2cmac_dat221,
                        ls2cmac_dat222,
                        ls2cmac_dat223,
                        ls2cmac_dat224,
                        ls2cmac_dat225,
                        ls2cmac_dat226,
                        ls2cmac_dat227,
                        ls2cmac_dat228,
                        ls2cmac_dat229,
                        ls2cmac_dat230,
                        ls2cmac_dat231,
                        ls2cmac_dat232,
                        ls2cmac_dat233,
                        ls2cmac_dat234,
                        ls2cmac_dat235,
                        ls2cmac_dat236,
                        ls2cmac_dat237,
                        ls2cmac_dat238,
                        ls2cmac_dat239,
                        ls2cmac_dat240,
                        ls2cmac_dat241,
                        ls2cmac_dat242,
                        ls2cmac_dat243,
                        ls2cmac_dat244,
                        ls2cmac_dat245,
                        ls2cmac_dat246,
                        ls2cmac_dat247,
                        ls2cmac_dat248,
                        ls2cmac_dat249,
                        ls2cmac_dat250,
                        ls2cmac_dat251,
                        ls2cmac_dat252,
                        ls2cmac_dat253,
                        ls2cmac_dat254,
                        ls2cmac_dat255,
                        ls2cmac_dat256,
                        ls2cmac_dat257,
                        ls2cmac_dat258,
                        ls2cmac_dat259,
                        ls2cmac_dat260,
                        ls2cmac_dat261,
                        ls2cmac_dat262,
                        ls2cmac_dat263,
                        ls2cmac_dat264,
                        ls2cmac_dat265,
                        ls2cmac_dat266,
                        ls2cmac_dat267,
                        ls2cmac_dat268,
                        ls2cmac_dat269,
                        ls2cmac_dat270,
                        ls2cmac_dat271,
                        ls2cmac_dat272,
                        ls2cmac_dat273,
                        ls2cmac_dat274,
                        ls2cmac_dat275,
                        ls2cmac_dat276,
                        ls2cmac_dat277,
                        ls2cmac_dat278,
                        ls2cmac_dat279,
                        ls2cmac_dat280,
                        ls2cmac_dat281,
                        ls2cmac_dat282,
                        ls2cmac_dat283,
                        ls2cmac_dat284,
                        ls2cmac_dat285,
                        ls2cmac_dat286,
                        ls2cmac_dat287,
                        ls2cmac_dat288,
                        ls2cmac_dat289,
                        ls2cmac_dat290,
                        ls2cmac_dat291,
                        ls2cmac_dat292,
                        ls2cmac_dat293,
                        ls2cmac_dat294,
                        ls2cmac_dat295,
                        ls2cmac_dat296,
                        ls2cmac_dat297,
                        ls2cmac_dat298,
                        ls2cmac_dat299,
                        ls2cmac_dat300,
                        ls2cmac_dat301,
                        ls2cmac_dat302,
                        ls2cmac_dat303,
                        ls2cmac_dat304,
                        ls2cmac_dat305,
                        ls2cmac_dat306,
                        ls2cmac_dat307,
                        ls2cmac_dat308,
                        ls2cmac_dat309,
                        ls2cmac_dat310,
                        ls2cmac_dat311,
                        ls2cmac_dat312,
                        ls2cmac_dat313,
                        ls2cmac_dat314,
                        ls2cmac_dat315,
                        ls2cmac_dat316,
                        ls2cmac_dat317,
                        ls2cmac_dat318,
                        ls2cmac_dat319,
                        ls2cmac_dat320,
                        ls2cmac_dat321,
                        ls2cmac_dat322,
                        ls2cmac_dat323,
                        ls2cmac_dat324,
                        ls2cmac_dat325,
                        ls2cmac_dat326,
                        ls2cmac_dat327,
                        ls2cmac_dat328,
                        ls2cmac_dat329,
                        ls2cmac_dat330,
                        ls2cmac_dat331,
                        ls2cmac_dat332,
                        ls2cmac_dat333,
                        ls2cmac_dat334,
                        ls2cmac_dat335,
                        ls2cmac_dat336,
                        ls2cmac_dat337,
                        ls2cmac_dat338,
                        ls2cmac_dat339,
                        ls2cmac_dat340,
                        ls2cmac_dat341,
                        ls2cmac_dat342,
                        ls2cmac_dat343,
                        ls2cmac_dat344,
                        ls2cmac_dat345,
                        ls2cmac_dat346,
                        ls2cmac_dat347,
                        ls2cmac_dat348,
                        ls2cmac_dat349,
                        ls2cmac_dat350,
                        ls2cmac_dat351,
                        ls2cmac_dat352,
                        ls2cmac_dat353,
                        ls2cmac_dat354,
                        ls2cmac_dat355,
                        ls2cmac_dat356,
                        ls2cmac_dat357,
                        ls2cmac_dat358,
                        ls2cmac_dat359,
                        ls2cmac_dat360,
                        ls2cmac_dat361,
                        ls2cmac_dat362,
                        ls2cmac_dat363,
                        ls2cmac_dat364,
                        ls2cmac_dat365,
                        ls2cmac_dat366,
                        ls2cmac_dat367,
                        ls2cmac_dat368,
                        ls2cmac_dat369,
                        ls2cmac_dat370,
                        ls2cmac_dat371,
                        ls2cmac_dat372,
                        ls2cmac_dat373,
                        ls2cmac_dat374,
                        ls2cmac_dat375,
                        ls2cmac_dat376,
                        ls2cmac_dat377,
                        ls2cmac_dat378,
                        ls2cmac_dat379,
                        ls2cmac_dat380,
                        ls2cmac_dat381,
                        ls2cmac_dat382,
                        ls2cmac_dat383,
                        ls2cmac_dat384,
                        ls2cmac_dat385,
                        ls2cmac_dat386,
                        ls2cmac_dat387,
                        ls2cmac_dat388,
                        ls2cmac_dat389,
                        ls2cmac_dat390,
                        ls2cmac_dat391,
                        ls2cmac_dat392,
                        ls2cmac_dat393,
                        ls2cmac_dat394,
                        ls2cmac_dat395,
                        ls2cmac_dat396,
                        ls2cmac_dat397,
                        ls2cmac_dat398,
                        ls2cmac_dat399,
                        ls2cmac_dat400,
                        ls2cmac_dat401,
                        ls2cmac_dat402,
                        ls2cmac_dat403,
                        ls2cmac_dat404,
                        ls2cmac_dat405,
                        ls2cmac_dat406,
                        ls2cmac_dat407,
                        ls2cmac_dat408,
                        ls2cmac_dat409,
                        ls2cmac_dat410,
                        ls2cmac_dat411,
                        ls2cmac_dat412,
                        ls2cmac_dat413,
                        ls2cmac_dat414,
                        ls2cmac_dat415,
                        ls2cmac_dat416,
                        ls2cmac_dat417,
                        ls2cmac_dat418,
                        ls2cmac_dat419,
                        ls2cmac_dat420,
                        ls2cmac_dat421,
                        ls2cmac_dat422,
                        ls2cmac_dat423,
                        ls2cmac_dat424,
                        ls2cmac_dat425,
                        ls2cmac_dat426,
                        ls2cmac_dat427,
                        ls2cmac_dat428,
                        ls2cmac_dat429,
                        ls2cmac_dat430,
                        ls2cmac_dat431,
                        ls2cmac_dat432,
                        ls2cmac_dat433,
                        ls2cmac_dat434,
                        ls2cmac_dat435,
                        ls2cmac_dat436,
                        ls2cmac_dat437,
                        ls2cmac_dat438,
                        ls2cmac_dat439,
                        ls2cmac_dat440,
                        ls2cmac_dat441,
                        ls2cmac_dat442,
                        ls2cmac_dat443,
                        ls2cmac_dat444,
                        ls2cmac_dat445,
                        ls2cmac_dat446,
                        ls2cmac_dat447,
                        ls2cmac_dat448,
                        ls2cmac_dat449,
                        ls2cmac_dat450,
                        ls2cmac_dat451,
                        ls2cmac_dat452,
                        ls2cmac_dat453,
                        ls2cmac_dat454,
                        ls2cmac_dat455,
                        ls2cmac_dat456,
                        ls2cmac_dat457,
                        ls2cmac_dat458,
                        ls2cmac_dat459,
                        ls2cmac_dat460,
                        ls2cmac_dat461,
                        ls2cmac_dat462,
                        ls2cmac_dat463,
                        ls2cmac_dat464,
                        ls2cmac_dat465,
                        ls2cmac_dat466,
                        ls2cmac_dat467,
                        ls2cmac_dat468,
                        ls2cmac_dat469,
                        ls2cmac_dat470,
                        ls2cmac_dat471,
                        ls2cmac_dat472,
                        ls2cmac_dat473,
                        ls2cmac_dat474,
                        ls2cmac_dat475,
                        ls2cmac_dat476,
                        ls2cmac_dat477,
                        ls2cmac_dat478,
                        ls2cmac_dat479,
                        ls2cmac_dat480,
                        ls2cmac_dat481,
                        ls2cmac_dat482,
                        ls2cmac_dat483,
                        ls2cmac_dat484,
                        ls2cmac_dat485,
                        ls2cmac_dat486,
                        ls2cmac_dat487,
                        ls2cmac_dat488,
                        ls2cmac_dat489,
                        ls2cmac_dat490,
                        ls2cmac_dat491,
                        ls2cmac_dat492,
                        ls2cmac_dat493,
                        ls2cmac_dat494,
                        ls2cmac_dat495,
                        ls2cmac_dat496,
                        ls2cmac_dat497,
                        ls2cmac_dat498,
                        ls2cmac_dat499,
                        ls2cmac_dat500,
                        ls2cmac_dat501,
                        ls2cmac_dat502,
                        ls2cmac_dat503,
                        ls2cmac_dat504,
                        ls2cmac_dat505,
                        ls2cmac_dat506,
                        ls2cmac_dat507,
                        ls2cmac_dat508,
                        ls2cmac_dat509,
                        ls2cmac_dat510,
                        ls2cmac_dat511,
                        ls2cmac_dat512,
                        ls2cmac_dat513,
                        ls2cmac_dat514,
                        ls2cmac_dat515,
                        ls2cmac_dat516,
                        ls2cmac_dat517,
                        ls2cmac_dat518,
                        ls2cmac_dat519,
                        ls2cmac_dat520,
                        ls2cmac_dat521,
                        ls2cmac_dat522,
                        ls2cmac_dat523,
                        ls2cmac_dat524,
                        ls2cmac_dat525,
                        ls2cmac_dat526,
                        ls2cmac_dat527,
                        ls2cmac_dat528,
                        ls2cmac_dat529,
                        ls2cmac_dat530,
                        ls2cmac_dat531,
                        ls2cmac_dat532,
                        ls2cmac_dat533,
                        ls2cmac_dat534,
                        ls2cmac_dat535,
                        ls2cmac_dat536,
                        ls2cmac_dat537,
                        ls2cmac_dat538,
                        ls2cmac_dat539,
                        ls2cmac_dat540,
                        ls2cmac_dat541,
                        ls2cmac_dat542,
                        ls2cmac_dat543,
                        ls2cmac_dat544,
                        ls2cmac_dat545,
                        ls2cmac_dat546,
                        ls2cmac_dat547,
                        ls2cmac_dat548,
                        ls2cmac_dat549,
                        ls2cmac_dat550,
                        ls2cmac_dat551,
                        ls2cmac_dat552,
                        ls2cmac_dat553,
                        ls2cmac_dat554,
                        ls2cmac_dat555,
                        ls2cmac_dat556,
                        ls2cmac_dat557,
                        ls2cmac_dat558,
                        ls2cmac_dat559,
                        ls2cmac_dat560,
                        ls2cmac_dat561,
                        ls2cmac_dat562,
                        ls2cmac_dat563,
                        ls2cmac_dat564,
                        ls2cmac_dat565,
                        ls2cmac_dat566,
                        ls2cmac_dat567,
                        ls2cmac_dat568,
                        ls2cmac_dat569,
                        ls2cmac_dat570,
                        ls2cmac_dat571,
                        ls2cmac_dat572,
                        ls2cmac_dat573,
                        ls2cmac_dat574,
                        ls2cmac_dat575,
                        ls2cmac_dat576,
                        ls2cmac_dat577,
                        ls2cmac_dat578,
                        ls2cmac_dat579,
                        ls2cmac_dat580,
                        ls2cmac_dat581,
                        ls2cmac_dat582,
                        ls2cmac_dat583,
                        ls2cmac_dat584,
                        ls2cmac_dat585,
                        ls2cmac_dat586,
                        ls2cmac_dat587,
                        ls2cmac_dat588,
                        ls2cmac_dat589,
                        ls2cmac_dat590,
                        ls2cmac_dat591,
                        ls2cmac_dat592,
                        ls2cmac_dat593,
                        ls2cmac_dat594,
                        ls2cmac_dat595,
                        ls2cmac_dat596,
                        ls2cmac_dat597,
                        ls2cmac_dat598,
                        ls2cmac_dat599,
                        ls2cmac_dat600,
                        ls2cmac_dat601,
                        ls2cmac_dat602,
                        ls2cmac_dat603,
                        ls2cmac_dat604,
                        ls2cmac_dat605,
                        ls2cmac_dat606,
                        ls2cmac_dat607,
                        ls2cmac_dat608,
                        ls2cmac_dat609,
                        ls2cmac_dat610,
                        ls2cmac_dat611,
                        ls2cmac_dat612,
                        ls2cmac_dat613,
                        ls2cmac_dat614,
                        ls2cmac_dat615,
                        ls2cmac_dat616,
                        ls2cmac_dat617,
                        ls2cmac_dat618,
                        ls2cmac_dat619,
                        ls2cmac_dat620,
                        ls2cmac_dat621,
                        ls2cmac_dat622,
                        ls2cmac_dat623,
                        ls2cmac_dat624,
                        ls2cmac_dat625,
                        ls2cmac_dat626,
                        ls2cmac_dat627,
                        ls2cmac_dat628,
                        ls2cmac_dat629,
                        ls2cmac_dat630,
                        ls2cmac_dat631,
                        ls2cmac_dat632,
                        ls2cmac_dat633,
                        ls2cmac_dat634,
                        ls2cmac_dat635,
                        ls2cmac_dat636,
                        ls2cmac_dat637,
                        ls2cmac_dat638,
                        ls2cmac_dat639,
                        ls2cmac_dat640,
                        ls2cmac_dat641,
                        ls2cmac_dat642,
                        ls2cmac_dat643,
                        ls2cmac_dat644,
                        ls2cmac_dat645,
                        ls2cmac_dat646,
                        ls2cmac_dat647,
                        ls2cmac_dat648,
                        ls2cmac_dat649,
                        ls2cmac_dat650,
                        ls2cmac_dat651,
                        ls2cmac_dat652,
                        ls2cmac_dat653,
                        ls2cmac_dat654,
                        ls2cmac_dat655,
                        ls2cmac_dat656,
                        ls2cmac_dat657,
                        ls2cmac_dat658,
                        ls2cmac_dat659,
                        ls2cmac_dat660,
                        ls2cmac_dat661,
                        ls2cmac_dat662,
                        ls2cmac_dat663,
                        ls2cmac_dat664,
                        ls2cmac_dat665,
                        ls2cmac_dat666,
                        ls2cmac_dat667,
                        ls2cmac_dat668,
                        ls2cmac_dat669,
                        ls2cmac_dat670,
                        ls2cmac_dat671,
                        ls2cmac_dat672,
                        ls2cmac_dat673,
                        ls2cmac_dat674,
                        ls2cmac_dat675,
                        ls2cmac_dat676,
                        ls2cmac_dat677,
                        ls2cmac_dat678,
                        ls2cmac_dat679,
                        ls2cmac_dat680,
                        ls2cmac_dat681,
                        ls2cmac_dat682,
                        ls2cmac_dat683,
                        ls2cmac_dat684,
                        ls2cmac_dat685,
                        ls2cmac_dat686,
                        ls2cmac_dat687,
                        ls2cmac_dat688,
                        ls2cmac_dat689,
                        ls2cmac_dat690,
                        ls2cmac_dat691,
                        ls2cmac_dat692,
                        ls2cmac_dat693,
                        ls2cmac_dat694,
                        ls2cmac_dat695,
                        ls2cmac_dat696,
                        ls2cmac_dat697,
                        ls2cmac_dat698,
                        ls2cmac_dat699,
                        ls2cmac_dat700,
                        ls2cmac_dat701,
                        ls2cmac_dat702,
                        ls2cmac_dat703,
                        ls2cmac_dat704,
                        ls2cmac_dat705,
                        ls2cmac_dat706,
                        ls2cmac_dat707,
                        ls2cmac_dat708,
                        ls2cmac_dat709,
                        ls2cmac_dat710,
                        ls2cmac_dat711,
                        ls2cmac_dat712,
                        ls2cmac_dat713,
                        ls2cmac_dat714,
                        ls2cmac_dat715,
                        ls2cmac_dat716,
                        ls2cmac_dat717,
                        ls2cmac_dat718,
                        ls2cmac_dat719,
                        ls2cmac_dat720,
                        ls2cmac_dat721,
                        ls2cmac_dat722,
                        ls2cmac_dat723,
                        ls2cmac_dat724,
                        ls2cmac_dat725,
                        ls2cmac_dat726,
                        ls2cmac_dat727,
                        ls2cmac_dat728,
                        ls2cmac_dat729,
                        ls2cmac_dat730,
                        ls2cmac_dat731,
                        ls2cmac_dat732,
                        ls2cmac_dat733,
                        ls2cmac_dat734,
                        ls2cmac_dat735,
                        ls2cmac_dat736,
                        ls2cmac_dat737,
                        ls2cmac_dat738,
                        ls2cmac_dat739,
                        ls2cmac_dat740,
                        ls2cmac_dat741,
                        ls2cmac_dat742,
                        ls2cmac_dat743,
                        ls2cmac_dat744,
                        ls2cmac_dat745,
                        ls2cmac_dat746,
                        ls2cmac_dat747,
                        ls2cmac_dat748,
                        ls2cmac_dat749,
                        ls2cmac_dat750,
                        ls2cmac_dat751,
                        ls2cmac_dat752,
                        ls2cmac_dat753,
                        ls2cmac_dat754,
                        ls2cmac_dat755,
                        ls2cmac_dat756,
                        ls2cmac_dat757,
                        ls2cmac_dat758,
                        ls2cmac_dat759,
                        ls2cmac_dat760,
                        ls2cmac_dat761,
                        ls2cmac_dat762,
                        ls2cmac_dat763,
                        ls2cmac_dat764,
                        ls2cmac_dat765,
                        ls2cmac_dat766,
                        ls2cmac_dat767,
                        ls2cmac_dat768,
                        ls2cmac_dat769,
                        ls2cmac_dat770,
                        ls2cmac_dat771,
                        ls2cmac_dat772,
                        ls2cmac_dat773,
                        ls2cmac_dat774,
                        ls2cmac_dat775,
                        ls2cmac_dat776,
                        ls2cmac_dat777,
                        ls2cmac_dat778,
                        ls2cmac_dat779,
                        ls2cmac_dat780,
                        ls2cmac_dat781,
                        ls2cmac_dat782,
                        ls2cmac_dat783,
                        ls2cmac_dat_size,
                        ls2cmac_wt0,
                        ls2cmac_wt1,
                        ls2cmac_wt2,
                        ls2cmac_wt3,
                        ls2cmac_wt4,
                        ls2cmac_wt5,
                        ls2cmac_wt6,
                        ls2cmac_wt7,
                        ls2cmac_wt8,
                        ls2cmac_wt9,
                        ls2cmac_wt10,
                        ls2cmac_wt11,
                        ls2cmac_wt12,
                        ls2cmac_wt13,
                        ls2cmac_wt14,
                        ls2cmac_wt15,
                        ls2cmac_wt16,
                        ls2cmac_wt17,
                        ls2cmac_wt18,
                        ls2cmac_wt19,
                        ls2cmac_wt20,
                        ls2cmac_wt21,
                        ls2cmac_wt22,
                        ls2cmac_wt23,
                        ls2cmac_wt24,
                        ls2cmac_wt_size,
                        conv2ls_output
                     );
    input       ytydla_core_clk;
    input       ytydla_core_rst_n;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat0;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat1;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat2;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat3;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat4;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat5;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat6;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat7;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat8;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat9;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat10;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat11;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat12;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat13;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat14;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat15;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat16;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat17;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat18;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat19;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat20;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat21;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat22;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat23;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat24;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat25;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat26;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat27;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat28;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat29;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat30;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat31;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat32;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat33;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat34;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat35;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat36;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat37;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat38;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat39;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat40;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat41;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat42;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat43;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat44;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat45;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat46;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat47;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat48;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat49;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat50;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat51;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat52;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat53;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat54;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat55;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat56;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat57;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat58;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat59;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat60;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat61;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat62;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat63;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat64;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat65;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat66;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat67;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat68;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat69;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat70;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat71;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat72;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat73;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat74;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat75;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat76;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat77;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat78;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat79;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat80;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat81;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat82;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat83;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat84;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat85;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat86;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat87;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat88;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat89;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat90;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat91;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat92;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat93;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat94;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat95;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat96;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat97;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat98;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat99;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat100;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat101;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat102;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat103;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat104;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat105;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat106;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat107;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat108;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat109;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat110;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat111;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat112;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat113;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat114;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat115;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat116;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat117;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat118;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat119;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat120;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat121;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat122;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat123;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat124;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat125;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat126;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat127;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat128;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat129;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat130;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat131;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat132;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat133;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat134;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat135;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat136;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat137;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat138;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat139;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat140;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat141;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat142;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat143;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat144;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat145;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat146;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat147;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat148;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat149;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat150;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat151;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat152;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat153;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat154;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat155;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat156;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat157;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat158;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat159;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat160;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat161;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat162;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat163;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat164;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat165;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat166;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat167;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat168;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat169;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat170;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat171;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat172;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat173;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat174;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat175;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat176;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat177;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat178;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat179;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat180;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat181;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat182;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat183;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat184;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat185;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat186;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat187;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat188;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat189;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat190;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat191;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat192;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat193;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat194;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat195;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat196;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat197;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat198;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat199;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat200;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat201;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat202;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat203;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat204;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat205;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat206;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat207;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat208;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat209;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat210;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat211;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat212;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat213;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat214;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat215;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat216;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat217;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat218;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat219;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat220;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat221;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat222;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat223;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat224;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat225;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat226;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat227;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat228;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat229;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat230;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat231;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat232;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat233;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat234;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat235;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat236;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat237;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat238;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat239;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat240;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat241;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat242;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat243;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat244;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat245;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat246;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat247;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat248;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat249;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat250;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat251;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat252;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat253;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat254;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat255;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat256;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat257;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat258;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat259;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat260;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat261;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat262;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat263;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat264;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat265;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat266;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat267;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat268;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat269;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat270;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat271;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat272;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat273;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat274;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat275;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat276;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat277;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat278;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat279;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat280;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat281;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat282;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat283;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat284;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat285;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat286;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat287;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat288;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat289;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat290;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat291;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat292;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat293;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat294;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat295;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat296;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat297;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat298;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat299;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat300;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat301;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat302;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat303;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat304;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat305;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat306;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat307;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat308;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat309;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat310;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat311;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat312;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat313;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat314;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat315;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat316;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat317;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat318;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat319;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat320;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat321;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat322;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat323;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat324;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat325;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat326;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat327;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat328;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat329;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat330;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat331;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat332;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat333;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat334;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat335;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat336;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat337;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat338;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat339;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat340;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat341;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat342;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat343;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat344;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat345;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat346;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat347;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat348;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat349;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat350;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat351;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat352;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat353;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat354;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat355;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat356;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat357;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat358;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat359;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat360;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat361;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat362;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat363;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat364;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat365;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat366;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat367;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat368;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat369;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat370;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat371;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat372;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat373;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat374;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat375;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat376;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat377;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat378;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat379;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat380;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat381;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat382;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat383;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat384;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat385;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat386;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat387;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat388;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat389;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat390;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat391;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat392;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat393;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat394;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat395;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat396;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat397;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat398;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat399;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat400;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat401;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat402;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat403;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat404;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat405;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat406;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat407;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat408;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat409;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat410;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat411;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat412;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat413;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat414;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat415;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat416;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat417;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat418;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat419;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat420;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat421;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat422;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat423;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat424;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat425;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat426;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat427;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat428;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat429;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat430;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat431;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat432;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat433;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat434;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat435;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat436;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat437;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat438;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat439;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat440;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat441;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat442;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat443;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat444;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat445;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat446;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat447;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat448;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat449;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat450;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat451;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat452;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat453;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat454;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat455;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat456;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat457;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat458;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat459;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat460;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat461;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat462;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat463;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat464;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat465;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat466;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat467;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat468;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat469;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat470;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat471;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat472;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat473;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat474;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat475;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat476;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat477;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat478;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat479;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat480;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat481;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat482;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat483;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat484;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat485;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat486;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat487;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat488;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat489;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat490;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat491;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat492;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat493;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat494;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat495;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat496;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat497;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat498;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat499;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat500;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat501;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat502;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat503;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat504;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat505;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat506;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat507;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat508;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat509;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat510;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat511;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat512;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat513;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat514;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat515;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat516;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat517;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat518;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat519;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat520;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat521;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat522;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat523;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat524;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat525;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat526;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat527;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat528;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat529;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat530;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat531;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat532;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat533;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat534;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat535;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat536;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat537;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat538;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat539;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat540;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat541;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat542;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat543;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat544;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat545;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat546;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat547;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat548;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat549;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat550;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat551;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat552;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat553;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat554;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat555;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat556;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat557;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat558;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat559;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat560;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat561;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat562;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat563;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat564;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat565;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat566;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat567;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat568;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat569;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat570;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat571;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat572;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat573;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat574;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat575;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat576;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat577;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat578;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat579;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat580;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat581;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat582;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat583;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat584;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat585;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat586;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat587;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat588;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat589;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat590;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat591;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat592;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat593;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat594;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat595;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat596;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat597;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat598;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat599;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat600;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat601;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat602;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat603;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat604;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat605;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat606;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat607;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat608;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat609;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat610;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat611;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat612;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat613;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat614;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat615;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat616;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat617;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat618;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat619;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat620;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat621;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat622;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat623;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat624;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat625;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat626;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat627;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat628;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat629;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat630;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat631;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat632;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat633;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat634;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat635;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat636;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat637;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat638;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat639;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat640;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat641;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat642;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat643;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat644;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat645;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat646;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat647;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat648;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat649;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat650;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat651;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat652;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat653;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat654;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat655;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat656;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat657;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat658;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat659;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat660;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat661;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat662;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat663;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat664;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat665;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat666;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat667;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat668;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat669;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat670;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat671;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat672;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat673;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat674;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat675;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat676;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat677;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat678;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat679;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat680;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat681;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat682;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat683;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat684;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat685;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat686;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat687;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat688;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat689;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat690;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat691;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat692;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat693;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat694;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat695;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat696;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat697;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat698;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat699;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat700;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat701;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat702;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat703;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat704;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat705;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat706;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat707;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat708;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat709;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat710;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat711;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat712;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat713;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat714;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat715;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat716;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat717;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat718;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat719;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat720;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat721;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat722;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat723;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat724;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat725;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat726;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat727;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat728;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat729;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat730;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat731;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat732;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat733;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat734;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat735;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat736;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat737;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat738;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat739;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat740;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat741;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat742;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat743;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat744;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat745;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat746;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat747;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat748;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat749;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat750;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat751;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat752;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat753;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat754;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat755;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat756;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat757;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat758;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat759;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat760;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat761;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat762;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat763;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat764;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat765;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat766;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat767;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat768;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat769;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat770;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat771;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat772;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat773;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat774;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat775;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat776;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat777;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat778;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat779;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat780;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat781;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat782;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_dat783;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt0;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt1;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt2;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt3;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt4;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt5;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt6;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt7;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt8;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt9;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt10;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt11;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt12;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt13;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt14;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt15;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt16;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt17;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt18;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt19;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt20;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt21;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt22;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt23;
    input    [YTYDLA_DATA_LENGTH - 1:0] ls2cmac_wt24;

        logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat0;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat1;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat2;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat3;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat4;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat5;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat6;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat7;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat8;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat9;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat10;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat11;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat12;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat13;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat14;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat15;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat16;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat17;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat18;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat19;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat20;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat21;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat22;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat23;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat24;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat25;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat26;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat27;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat28;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat29;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat30;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat31;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat32;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat33;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat34;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat35;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat36;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat37;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat38;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat39;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat40;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat41;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat42;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat43;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat44;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat45;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat46;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat47;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat48;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat49;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat50;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat51;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat52;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat53;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat54;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat55;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat56;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat57;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat58;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat59;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat60;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat61;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat62;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat63;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat64;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat65;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat66;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat67;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat68;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat69;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat70;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat71;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat72;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat73;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat74;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat75;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat76;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat77;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat78;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat79;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat80;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat81;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat82;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat83;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat84;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat85;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat86;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat87;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat88;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat89;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat90;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat91;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat92;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat93;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat94;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat95;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat96;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat97;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat98;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat99;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat100;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat101;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat102;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat103;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat104;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat105;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat106;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat107;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat108;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat109;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat110;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat111;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat112;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat113;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat114;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat115;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat116;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat117;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat118;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat119;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat120;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat121;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat122;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat123;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat124;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat125;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat126;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat127;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat128;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat129;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat130;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat131;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat132;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat133;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat134;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat135;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat136;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat137;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat138;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat139;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat140;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat141;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat142;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat143;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat144;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat145;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat146;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat147;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat148;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat149;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat150;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat151;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat152;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat153;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat154;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat155;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat156;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat157;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat158;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat159;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat160;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat161;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat162;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat163;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat164;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat165;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat166;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat167;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat168;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat169;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat170;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat171;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat172;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat173;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat174;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat175;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat176;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat177;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat178;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat179;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat180;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat181;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat182;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat183;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat184;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat185;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat186;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat187;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat188;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat189;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat190;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat191;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat192;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat193;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat194;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat195;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat196;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat197;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat198;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat199;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat200;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat201;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat202;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat203;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat204;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat205;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat206;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat207;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat208;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat209;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat210;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat211;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat212;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat213;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat214;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat215;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat216;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat217;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat218;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat219;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat220;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat221;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat222;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat223;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat224;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat225;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat226;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat227;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat228;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat229;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat230;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat231;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat232;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat233;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat234;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat235;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat236;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat237;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat238;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat239;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat240;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat241;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat242;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat243;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat244;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat245;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat246;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat247;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat248;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat249;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat250;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat251;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat252;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat253;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat254;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat255;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat256;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat257;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat258;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat259;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat260;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat261;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat262;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat263;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat264;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat265;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat266;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat267;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat268;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat269;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat270;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat271;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat272;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat273;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat274;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat275;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat276;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat277;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat278;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat279;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat280;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat281;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat282;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat283;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat284;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat285;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat286;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat287;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat288;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat289;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat290;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat291;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat292;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat293;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat294;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat295;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat296;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat297;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat298;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat299;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat300;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat301;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat302;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat303;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat304;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat305;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat306;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat307;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat308;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat309;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat310;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat311;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat312;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat313;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat314;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat315;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat316;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat317;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat318;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat319;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat320;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat321;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat322;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat323;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat324;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat325;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat326;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat327;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat328;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat329;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat330;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat331;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat332;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat333;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat334;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat335;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat336;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat337;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat338;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat339;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat340;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat341;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat342;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat343;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat344;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat345;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat346;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat347;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat348;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat349;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat350;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat351;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat352;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat353;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat354;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat355;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat356;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat357;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat358;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat359;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat360;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat361;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat362;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat363;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat364;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat365;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat366;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat367;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat368;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat369;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat370;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat371;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat372;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat373;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat374;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat375;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat376;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat377;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat378;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat379;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat380;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat381;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat382;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat383;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat384;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat385;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat386;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat387;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat388;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat389;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat390;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat391;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat392;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat393;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat394;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat395;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat396;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat397;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat398;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat399;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat400;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat401;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat402;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat403;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat404;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat405;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat406;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat407;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat408;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat409;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat410;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat411;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat412;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat413;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat414;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat415;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat416;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat417;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat418;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat419;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat420;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat421;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat422;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat423;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat424;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat425;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat426;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat427;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat428;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat429;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat430;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat431;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat432;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat433;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat434;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat435;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat436;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat437;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat438;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat439;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat440;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat441;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat442;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat443;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat444;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat445;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat446;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat447;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat448;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat449;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat450;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat451;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat452;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat453;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat454;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat455;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat456;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat457;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat458;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat459;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat460;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat461;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat462;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat463;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat464;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat465;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat466;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat467;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat468;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat469;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat470;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat471;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat472;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat473;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat474;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat475;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat476;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat477;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat478;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat479;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat480;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat481;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat482;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat483;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat484;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat485;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat486;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat487;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat488;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat489;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat490;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat491;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat492;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat493;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat494;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat495;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat496;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat497;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat498;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat499;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat500;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat501;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat502;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat503;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat504;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat505;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat506;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat507;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat508;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat509;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat510;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat511;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat512;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat513;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat514;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat515;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat516;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat517;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat518;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat519;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat520;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat521;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat522;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat523;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat524;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat525;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat526;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat527;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat528;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat529;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat530;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat531;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat532;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat533;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat534;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat535;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat536;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat537;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat538;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat539;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat540;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat541;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat542;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat543;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat544;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat545;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat546;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat547;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat548;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat549;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat550;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat551;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat552;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat553;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat554;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat555;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat556;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat557;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat558;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat559;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat560;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat561;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat562;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat563;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat564;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat565;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat566;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat567;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat568;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat569;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat570;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat571;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat572;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat573;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat574;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat575;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat576;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat577;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat578;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat579;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat580;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat581;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat582;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat583;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat584;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat585;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat586;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat587;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat588;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat589;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat590;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat591;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat592;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat593;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat594;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat595;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat596;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat597;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat598;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat599;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat600;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat601;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat602;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat603;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat604;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat605;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat606;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat607;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat608;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat609;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat610;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat611;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat612;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat613;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat614;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat615;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat616;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat617;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat618;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat619;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat620;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat621;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat622;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat623;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat624;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat625;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat626;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat627;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat628;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat629;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat630;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat631;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat632;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat633;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat634;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat635;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat636;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat637;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat638;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat639;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat640;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat641;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat642;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat643;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat644;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat645;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat646;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat647;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat648;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat649;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat650;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat651;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat652;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat653;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat654;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat655;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat656;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat657;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat658;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat659;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat660;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat661;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat662;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat663;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat664;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat665;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat666;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat667;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat668;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat669;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat670;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat671;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat672;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat673;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat674;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat675;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat676;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat677;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat678;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat679;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat680;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat681;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat682;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat683;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat684;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat685;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat686;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat687;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat688;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat689;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat690;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat691;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat692;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat693;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat694;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat695;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat696;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat697;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat698;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat699;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat700;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat701;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat702;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat703;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat704;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat705;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat706;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat707;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat708;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat709;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat710;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat711;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat712;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat713;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat714;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat715;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat716;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat717;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat718;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat719;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat720;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat721;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat722;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat723;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat724;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat725;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat726;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat727;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat728;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat729;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat730;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat731;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat732;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat733;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat734;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat735;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat736;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat737;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat738;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat739;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat740;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat741;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat742;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat743;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat744;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat745;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat746;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat747;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat748;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat749;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat750;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat751;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat752;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat753;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat754;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat755;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat756;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat757;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat758;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat759;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat760;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat761;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat762;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat763;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat764;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat765;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat766;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat767;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat768;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat769;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat770;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat771;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat772;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat773;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat774;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat775;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat776;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat777;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat778;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat779;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat780;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat781;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat782;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_dat783;

    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt0;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt1;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt2;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt3;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt4;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt5;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt6;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt7;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt8;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt9;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt10;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt11;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt12;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt13;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt14;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt15;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt16;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt17;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt18;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt19;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt20;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt21;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt22;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt23;
    logic    [YTYDLA_DATA_LENGTH - 1:0] conv_wt24;

    logic      [24:0]                   conv2cmac_dat_bigmap;
    logic      [24:0]                   conv2cmac_wt_bitmap;

    assign      conv2cmac_dat_bigmap = 25'1ffffff;
    assign      conv2cmac_wt_bitmap = 25'1ffffff;

    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt0 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt0 <= ls2cmac_wt0;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt1 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt1 <= ls2cmac_wt1;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt2 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt2 <= ls2cmac_wt2;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt3 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt3 <= ls2cmac_wt3;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt4 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt4 <= ls2cmac_wt4;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt5 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt5 <= ls2cmac_wt5;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt6 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt6 <= ls2cmac_wt6;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt7 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt7 <= ls2cmac_wt7;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt8 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt8 <= ls2cmac_wt8;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt9 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt9 <= ls2cmac_wt9;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt10 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt10 <= ls2cmac_wt10;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt11 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt11 <= ls2cmac_wt11;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt12 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt12 <= ls2cmac_wt12;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt13 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt13 <= ls2cmac_wt13;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt14 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt14 <= ls2cmac_wt14;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt15 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt15 <= ls2cmac_wt15;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt16 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt16 <= ls2cmac_wt16;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt17 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt17 <= ls2cmac_wt17;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt18 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt18 <= ls2cmac_wt18;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt19 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt19 <= ls2cmac_wt19;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt20 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt20 <= ls2cmac_wt20;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt21 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt21 <= ls2cmac_wt21;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt22 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt22 <= ls2cmac_wt22;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt23 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt23 <= ls2cmac_wt23;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_wt24 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_wt24 <= ls2cmac_wt24;
        end
    end

        always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat0 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat0 <= ls2cmac_dat0;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat1 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat1 <= ls2cmac_dat1;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat2 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat2 <= ls2cmac_dat2;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat3 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat3 <= ls2cmac_dat3;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat4 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat4 <= ls2cmac_dat4;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat5 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat5 <= ls2cmac_dat5;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat6 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat6 <= ls2cmac_dat6;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat7 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat7 <= ls2cmac_dat7;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat8 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat8 <= ls2cmac_dat8;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat9 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat9 <= ls2cmac_dat9;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat10 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat10 <= ls2cmac_dat10;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat11 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat11 <= ls2cmac_dat11;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat12 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat12 <= ls2cmac_dat12;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat13 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat13 <= ls2cmac_dat13;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat14 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat14 <= ls2cmac_dat14;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat15 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat15 <= ls2cmac_dat15;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat16 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat16 <= ls2cmac_dat16;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat17 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat17 <= ls2cmac_dat17;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat18 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat18 <= ls2cmac_dat18;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat19 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat19 <= ls2cmac_dat19;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat20 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat20 <= ls2cmac_dat20;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat21 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat21 <= ls2cmac_dat21;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat22 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat22 <= ls2cmac_dat22;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat23 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat23 <= ls2cmac_dat23;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat24 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat24 <= ls2cmac_dat24;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat25 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat25 <= ls2cmac_dat25;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat26 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat26 <= ls2cmac_dat26;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat27 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat27 <= ls2cmac_dat27;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat28 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat28 <= ls2cmac_dat28;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat29 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat29 <= ls2cmac_dat29;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat30 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat30 <= ls2cmac_dat30;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat31 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat31 <= ls2cmac_dat31;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat32 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat32 <= ls2cmac_dat32;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat33 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat33 <= ls2cmac_dat33;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat34 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat34 <= ls2cmac_dat34;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat35 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat35 <= ls2cmac_dat35;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat36 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat36 <= ls2cmac_dat36;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat37 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat37 <= ls2cmac_dat37;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat38 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat38 <= ls2cmac_dat38;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat39 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat39 <= ls2cmac_dat39;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat40 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat40 <= ls2cmac_dat40;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat41 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat41 <= ls2cmac_dat41;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat42 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat42 <= ls2cmac_dat42;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat43 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat43 <= ls2cmac_dat43;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat44 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat44 <= ls2cmac_dat44;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat45 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat45 <= ls2cmac_dat45;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat46 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat46 <= ls2cmac_dat46;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat47 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat47 <= ls2cmac_dat47;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat48 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat48 <= ls2cmac_dat48;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat49 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat49 <= ls2cmac_dat49;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat50 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat50 <= ls2cmac_dat50;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat51 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat51 <= ls2cmac_dat51;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat52 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat52 <= ls2cmac_dat52;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat53 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat53 <= ls2cmac_dat53;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat54 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat54 <= ls2cmac_dat54;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat55 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat55 <= ls2cmac_dat55;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat56 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat56 <= ls2cmac_dat56;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat57 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat57 <= ls2cmac_dat57;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat58 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat58 <= ls2cmac_dat58;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat59 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat59 <= ls2cmac_dat59;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat60 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat60 <= ls2cmac_dat60;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat61 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat61 <= ls2cmac_dat61;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat62 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat62 <= ls2cmac_dat62;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat63 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat63 <= ls2cmac_dat63;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat64 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat64 <= ls2cmac_dat64;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat65 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat65 <= ls2cmac_dat65;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat66 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat66 <= ls2cmac_dat66;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat67 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat67 <= ls2cmac_dat67;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat68 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat68 <= ls2cmac_dat68;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat69 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat69 <= ls2cmac_dat69;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat70 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat70 <= ls2cmac_dat70;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat71 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat71 <= ls2cmac_dat71;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat72 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat72 <= ls2cmac_dat72;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat73 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat73 <= ls2cmac_dat73;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat74 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat74 <= ls2cmac_dat74;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat75 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat75 <= ls2cmac_dat75;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat76 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat76 <= ls2cmac_dat76;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat77 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat77 <= ls2cmac_dat77;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat78 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat78 <= ls2cmac_dat78;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat79 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat79 <= ls2cmac_dat79;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat80 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat80 <= ls2cmac_dat80;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat81 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat81 <= ls2cmac_dat81;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat82 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat82 <= ls2cmac_dat82;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat83 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat83 <= ls2cmac_dat83;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat84 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat84 <= ls2cmac_dat84;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat85 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat85 <= ls2cmac_dat85;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat86 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat86 <= ls2cmac_dat86;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat87 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat87 <= ls2cmac_dat87;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat88 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat88 <= ls2cmac_dat88;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat89 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat89 <= ls2cmac_dat89;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat90 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat90 <= ls2cmac_dat90;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat91 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat91 <= ls2cmac_dat91;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat92 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat92 <= ls2cmac_dat92;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat93 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat93 <= ls2cmac_dat93;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat94 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat94 <= ls2cmac_dat94;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat95 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat95 <= ls2cmac_dat95;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat96 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat96 <= ls2cmac_dat96;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat97 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat97 <= ls2cmac_dat97;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat98 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat98 <= ls2cmac_dat98;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat99 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat99 <= ls2cmac_dat99;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat100 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat100 <= ls2cmac_dat100;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat101 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat101 <= ls2cmac_dat101;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat102 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat102 <= ls2cmac_dat102;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat103 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat103 <= ls2cmac_dat103;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat104 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat104 <= ls2cmac_dat104;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat105 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat105 <= ls2cmac_dat105;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat106 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat106 <= ls2cmac_dat106;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat107 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat107 <= ls2cmac_dat107;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat108 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat108 <= ls2cmac_dat108;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat109 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat109 <= ls2cmac_dat109;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat110 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat110 <= ls2cmac_dat110;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat111 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat111 <= ls2cmac_dat111;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat112 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat112 <= ls2cmac_dat112;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat113 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat113 <= ls2cmac_dat113;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat114 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat114 <= ls2cmac_dat114;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat115 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat115 <= ls2cmac_dat115;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat116 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat116 <= ls2cmac_dat116;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat117 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat117 <= ls2cmac_dat117;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat118 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat118 <= ls2cmac_dat118;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat119 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat119 <= ls2cmac_dat119;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat120 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat120 <= ls2cmac_dat120;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat121 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat121 <= ls2cmac_dat121;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat122 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat122 <= ls2cmac_dat122;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat123 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat123 <= ls2cmac_dat123;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat124 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat124 <= ls2cmac_dat124;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat125 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat125 <= ls2cmac_dat125;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat126 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat126 <= ls2cmac_dat126;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat127 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat127 <= ls2cmac_dat127;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat128 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat128 <= ls2cmac_dat128;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat129 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat129 <= ls2cmac_dat129;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat130 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat130 <= ls2cmac_dat130;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat131 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat131 <= ls2cmac_dat131;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat132 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat132 <= ls2cmac_dat132;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat133 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat133 <= ls2cmac_dat133;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat134 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat134 <= ls2cmac_dat134;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat135 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat135 <= ls2cmac_dat135;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat136 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat136 <= ls2cmac_dat136;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat137 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat137 <= ls2cmac_dat137;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat138 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat138 <= ls2cmac_dat138;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat139 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat139 <= ls2cmac_dat139;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat140 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat140 <= ls2cmac_dat140;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat141 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat141 <= ls2cmac_dat141;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat142 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat142 <= ls2cmac_dat142;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat143 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat143 <= ls2cmac_dat143;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat144 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat144 <= ls2cmac_dat144;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat145 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat145 <= ls2cmac_dat145;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat146 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat146 <= ls2cmac_dat146;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat147 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat147 <= ls2cmac_dat147;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat148 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat148 <= ls2cmac_dat148;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat149 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat149 <= ls2cmac_dat149;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat150 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat150 <= ls2cmac_dat150;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat151 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat151 <= ls2cmac_dat151;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat152 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat152 <= ls2cmac_dat152;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat153 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat153 <= ls2cmac_dat153;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat154 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat154 <= ls2cmac_dat154;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat155 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat155 <= ls2cmac_dat155;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat156 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat156 <= ls2cmac_dat156;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat157 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat157 <= ls2cmac_dat157;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat158 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat158 <= ls2cmac_dat158;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat159 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat159 <= ls2cmac_dat159;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat160 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat160 <= ls2cmac_dat160;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat161 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat161 <= ls2cmac_dat161;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat162 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat162 <= ls2cmac_dat162;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat163 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat163 <= ls2cmac_dat163;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat164 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat164 <= ls2cmac_dat164;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat165 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat165 <= ls2cmac_dat165;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat166 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat166 <= ls2cmac_dat166;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat167 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat167 <= ls2cmac_dat167;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat168 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat168 <= ls2cmac_dat168;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat169 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat169 <= ls2cmac_dat169;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat170 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat170 <= ls2cmac_dat170;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat171 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat171 <= ls2cmac_dat171;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat172 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat172 <= ls2cmac_dat172;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat173 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat173 <= ls2cmac_dat173;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat174 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat174 <= ls2cmac_dat174;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat175 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat175 <= ls2cmac_dat175;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat176 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat176 <= ls2cmac_dat176;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat177 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat177 <= ls2cmac_dat177;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat178 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat178 <= ls2cmac_dat178;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat179 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat179 <= ls2cmac_dat179;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat180 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat180 <= ls2cmac_dat180;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat181 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat181 <= ls2cmac_dat181;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat182 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat182 <= ls2cmac_dat182;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat183 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat183 <= ls2cmac_dat183;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat184 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat184 <= ls2cmac_dat184;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat185 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat185 <= ls2cmac_dat185;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat186 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat186 <= ls2cmac_dat186;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat187 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat187 <= ls2cmac_dat187;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat188 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat188 <= ls2cmac_dat188;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat189 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat189 <= ls2cmac_dat189;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat190 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat190 <= ls2cmac_dat190;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat191 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat191 <= ls2cmac_dat191;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat192 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat192 <= ls2cmac_dat192;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat193 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat193 <= ls2cmac_dat193;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat194 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat194 <= ls2cmac_dat194;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat195 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat195 <= ls2cmac_dat195;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat196 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat196 <= ls2cmac_dat196;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat197 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat197 <= ls2cmac_dat197;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat198 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat198 <= ls2cmac_dat198;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat199 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat199 <= ls2cmac_dat199;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat200 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat200 <= ls2cmac_dat200;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat201 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat201 <= ls2cmac_dat201;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat202 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat202 <= ls2cmac_dat202;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat203 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat203 <= ls2cmac_dat203;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat204 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat204 <= ls2cmac_dat204;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat205 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat205 <= ls2cmac_dat205;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat206 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat206 <= ls2cmac_dat206;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat207 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat207 <= ls2cmac_dat207;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat208 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat208 <= ls2cmac_dat208;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat209 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat209 <= ls2cmac_dat209;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat210 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat210 <= ls2cmac_dat210;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat211 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat211 <= ls2cmac_dat211;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat212 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat212 <= ls2cmac_dat212;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat213 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat213 <= ls2cmac_dat213;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat214 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat214 <= ls2cmac_dat214;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat215 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat215 <= ls2cmac_dat215;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat216 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat216 <= ls2cmac_dat216;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat217 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat217 <= ls2cmac_dat217;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat218 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat218 <= ls2cmac_dat218;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat219 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat219 <= ls2cmac_dat219;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat220 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat220 <= ls2cmac_dat220;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat221 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat221 <= ls2cmac_dat221;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat222 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat222 <= ls2cmac_dat222;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat223 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat223 <= ls2cmac_dat223;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat224 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat224 <= ls2cmac_dat224;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat225 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat225 <= ls2cmac_dat225;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat226 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat226 <= ls2cmac_dat226;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat227 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat227 <= ls2cmac_dat227;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat228 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat228 <= ls2cmac_dat228;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat229 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat229 <= ls2cmac_dat229;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat230 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat230 <= ls2cmac_dat230;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat231 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat231 <= ls2cmac_dat231;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat232 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat232 <= ls2cmac_dat232;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat233 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat233 <= ls2cmac_dat233;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat234 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat234 <= ls2cmac_dat234;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat235 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat235 <= ls2cmac_dat235;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat236 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat236 <= ls2cmac_dat236;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat237 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat237 <= ls2cmac_dat237;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat238 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat238 <= ls2cmac_dat238;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat239 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat239 <= ls2cmac_dat239;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat240 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat240 <= ls2cmac_dat240;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat241 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat241 <= ls2cmac_dat241;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat242 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat242 <= ls2cmac_dat242;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat243 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat243 <= ls2cmac_dat243;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat244 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat244 <= ls2cmac_dat244;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat245 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat245 <= ls2cmac_dat245;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat246 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat246 <= ls2cmac_dat246;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat247 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat247 <= ls2cmac_dat247;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat248 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat248 <= ls2cmac_dat248;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat249 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat249 <= ls2cmac_dat249;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat250 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat250 <= ls2cmac_dat250;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat251 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat251 <= ls2cmac_dat251;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat252 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat252 <= ls2cmac_dat252;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat253 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat253 <= ls2cmac_dat253;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat254 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat254 <= ls2cmac_dat254;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat255 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat255 <= ls2cmac_dat255;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat256 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat256 <= ls2cmac_dat256;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat257 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat257 <= ls2cmac_dat257;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat258 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat258 <= ls2cmac_dat258;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat259 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat259 <= ls2cmac_dat259;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat260 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat260 <= ls2cmac_dat260;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat261 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat261 <= ls2cmac_dat261;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat262 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat262 <= ls2cmac_dat262;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat263 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat263 <= ls2cmac_dat263;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat264 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat264 <= ls2cmac_dat264;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat265 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat265 <= ls2cmac_dat265;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat266 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat266 <= ls2cmac_dat266;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat267 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat267 <= ls2cmac_dat267;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat268 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat268 <= ls2cmac_dat268;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat269 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat269 <= ls2cmac_dat269;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat270 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat270 <= ls2cmac_dat270;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat271 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat271 <= ls2cmac_dat271;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat272 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat272 <= ls2cmac_dat272;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat273 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat273 <= ls2cmac_dat273;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat274 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat274 <= ls2cmac_dat274;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat275 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat275 <= ls2cmac_dat275;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat276 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat276 <= ls2cmac_dat276;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat277 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat277 <= ls2cmac_dat277;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat278 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat278 <= ls2cmac_dat278;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat279 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat279 <= ls2cmac_dat279;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat280 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat280 <= ls2cmac_dat280;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat281 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat281 <= ls2cmac_dat281;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat282 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat282 <= ls2cmac_dat282;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat283 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat283 <= ls2cmac_dat283;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat284 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat284 <= ls2cmac_dat284;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat285 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat285 <= ls2cmac_dat285;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat286 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat286 <= ls2cmac_dat286;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat287 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat287 <= ls2cmac_dat287;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat288 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat288 <= ls2cmac_dat288;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat289 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat289 <= ls2cmac_dat289;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat290 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat290 <= ls2cmac_dat290;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat291 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat291 <= ls2cmac_dat291;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat292 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat292 <= ls2cmac_dat292;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat293 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat293 <= ls2cmac_dat293;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat294 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat294 <= ls2cmac_dat294;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat295 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat295 <= ls2cmac_dat295;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat296 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat296 <= ls2cmac_dat296;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat297 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat297 <= ls2cmac_dat297;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat298 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat298 <= ls2cmac_dat298;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat299 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat299 <= ls2cmac_dat299;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat300 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat300 <= ls2cmac_dat300;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat301 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat301 <= ls2cmac_dat301;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat302 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat302 <= ls2cmac_dat302;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat303 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat303 <= ls2cmac_dat303;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat304 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat304 <= ls2cmac_dat304;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat305 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat305 <= ls2cmac_dat305;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat306 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat306 <= ls2cmac_dat306;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat307 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat307 <= ls2cmac_dat307;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat308 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat308 <= ls2cmac_dat308;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat309 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat309 <= ls2cmac_dat309;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat310 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat310 <= ls2cmac_dat310;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat311 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat311 <= ls2cmac_dat311;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat312 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat312 <= ls2cmac_dat312;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat313 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat313 <= ls2cmac_dat313;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat314 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat314 <= ls2cmac_dat314;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat315 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat315 <= ls2cmac_dat315;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat316 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat316 <= ls2cmac_dat316;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat317 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat317 <= ls2cmac_dat317;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat318 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat318 <= ls2cmac_dat318;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat319 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat319 <= ls2cmac_dat319;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat320 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat320 <= ls2cmac_dat320;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat321 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat321 <= ls2cmac_dat321;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat322 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat322 <= ls2cmac_dat322;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat323 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat323 <= ls2cmac_dat323;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat324 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat324 <= ls2cmac_dat324;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat325 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat325 <= ls2cmac_dat325;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat326 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat326 <= ls2cmac_dat326;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat327 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat327 <= ls2cmac_dat327;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat328 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat328 <= ls2cmac_dat328;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat329 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat329 <= ls2cmac_dat329;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat330 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat330 <= ls2cmac_dat330;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat331 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat331 <= ls2cmac_dat331;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat332 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat332 <= ls2cmac_dat332;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat333 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat333 <= ls2cmac_dat333;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat334 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat334 <= ls2cmac_dat334;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat335 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat335 <= ls2cmac_dat335;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat336 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat336 <= ls2cmac_dat336;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat337 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat337 <= ls2cmac_dat337;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat338 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat338 <= ls2cmac_dat338;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat339 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat339 <= ls2cmac_dat339;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat340 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat340 <= ls2cmac_dat340;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat341 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat341 <= ls2cmac_dat341;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat342 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat342 <= ls2cmac_dat342;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat343 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat343 <= ls2cmac_dat343;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat344 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat344 <= ls2cmac_dat344;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat345 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat345 <= ls2cmac_dat345;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat346 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat346 <= ls2cmac_dat346;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat347 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat347 <= ls2cmac_dat347;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat348 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat348 <= ls2cmac_dat348;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat349 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat349 <= ls2cmac_dat349;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat350 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat350 <= ls2cmac_dat350;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat351 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat351 <= ls2cmac_dat351;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat352 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat352 <= ls2cmac_dat352;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat353 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat353 <= ls2cmac_dat353;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat354 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat354 <= ls2cmac_dat354;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat355 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat355 <= ls2cmac_dat355;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat356 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat356 <= ls2cmac_dat356;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat357 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat357 <= ls2cmac_dat357;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat358 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat358 <= ls2cmac_dat358;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat359 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat359 <= ls2cmac_dat359;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat360 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat360 <= ls2cmac_dat360;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat361 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat361 <= ls2cmac_dat361;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat362 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat362 <= ls2cmac_dat362;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat363 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat363 <= ls2cmac_dat363;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat364 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat364 <= ls2cmac_dat364;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat365 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat365 <= ls2cmac_dat365;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat366 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat366 <= ls2cmac_dat366;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat367 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat367 <= ls2cmac_dat367;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat368 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat368 <= ls2cmac_dat368;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat369 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat369 <= ls2cmac_dat369;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat370 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat370 <= ls2cmac_dat370;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat371 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat371 <= ls2cmac_dat371;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat372 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat372 <= ls2cmac_dat372;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat373 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat373 <= ls2cmac_dat373;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat374 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat374 <= ls2cmac_dat374;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat375 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat375 <= ls2cmac_dat375;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat376 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat376 <= ls2cmac_dat376;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat377 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat377 <= ls2cmac_dat377;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat378 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat378 <= ls2cmac_dat378;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat379 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat379 <= ls2cmac_dat379;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat380 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat380 <= ls2cmac_dat380;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat381 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat381 <= ls2cmac_dat381;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat382 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat382 <= ls2cmac_dat382;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat383 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat383 <= ls2cmac_dat383;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat384 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat384 <= ls2cmac_dat384;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat385 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat385 <= ls2cmac_dat385;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat386 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat386 <= ls2cmac_dat386;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat387 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat387 <= ls2cmac_dat387;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat388 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat388 <= ls2cmac_dat388;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat389 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat389 <= ls2cmac_dat389;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat390 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat390 <= ls2cmac_dat390;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat391 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat391 <= ls2cmac_dat391;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat392 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat392 <= ls2cmac_dat392;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat393 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat393 <= ls2cmac_dat393;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat394 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat394 <= ls2cmac_dat394;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat395 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat395 <= ls2cmac_dat395;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat396 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat396 <= ls2cmac_dat396;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat397 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat397 <= ls2cmac_dat397;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat398 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat398 <= ls2cmac_dat398;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat399 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat399 <= ls2cmac_dat399;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat400 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat400 <= ls2cmac_dat400;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat401 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat401 <= ls2cmac_dat401;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat402 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat402 <= ls2cmac_dat402;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat403 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat403 <= ls2cmac_dat403;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat404 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat404 <= ls2cmac_dat404;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat405 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat405 <= ls2cmac_dat405;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat406 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat406 <= ls2cmac_dat406;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat407 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat407 <= ls2cmac_dat407;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat408 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat408 <= ls2cmac_dat408;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat409 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat409 <= ls2cmac_dat409;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat410 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat410 <= ls2cmac_dat410;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat411 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat411 <= ls2cmac_dat411;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat412 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat412 <= ls2cmac_dat412;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat413 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat413 <= ls2cmac_dat413;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat414 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat414 <= ls2cmac_dat414;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat415 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat415 <= ls2cmac_dat415;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat416 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat416 <= ls2cmac_dat416;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat417 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat417 <= ls2cmac_dat417;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat418 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat418 <= ls2cmac_dat418;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat419 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat419 <= ls2cmac_dat419;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat420 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat420 <= ls2cmac_dat420;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat421 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat421 <= ls2cmac_dat421;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat422 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat422 <= ls2cmac_dat422;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat423 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat423 <= ls2cmac_dat423;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat424 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat424 <= ls2cmac_dat424;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat425 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat425 <= ls2cmac_dat425;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat426 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat426 <= ls2cmac_dat426;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat427 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat427 <= ls2cmac_dat427;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat428 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat428 <= ls2cmac_dat428;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat429 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat429 <= ls2cmac_dat429;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat430 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat430 <= ls2cmac_dat430;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat431 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat431 <= ls2cmac_dat431;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat432 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat432 <= ls2cmac_dat432;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat433 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat433 <= ls2cmac_dat433;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat434 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat434 <= ls2cmac_dat434;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat435 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat435 <= ls2cmac_dat435;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat436 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat436 <= ls2cmac_dat436;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat437 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat437 <= ls2cmac_dat437;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat438 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat438 <= ls2cmac_dat438;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat439 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat439 <= ls2cmac_dat439;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat440 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat440 <= ls2cmac_dat440;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat441 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat441 <= ls2cmac_dat441;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat442 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat442 <= ls2cmac_dat442;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat443 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat443 <= ls2cmac_dat443;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat444 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat444 <= ls2cmac_dat444;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat445 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat445 <= ls2cmac_dat445;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat446 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat446 <= ls2cmac_dat446;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat447 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat447 <= ls2cmac_dat447;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat448 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat448 <= ls2cmac_dat448;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat449 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat449 <= ls2cmac_dat449;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat450 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat450 <= ls2cmac_dat450;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat451 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat451 <= ls2cmac_dat451;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat452 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat452 <= ls2cmac_dat452;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat453 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat453 <= ls2cmac_dat453;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat454 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat454 <= ls2cmac_dat454;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat455 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat455 <= ls2cmac_dat455;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat456 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat456 <= ls2cmac_dat456;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat457 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat457 <= ls2cmac_dat457;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat458 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat458 <= ls2cmac_dat458;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat459 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat459 <= ls2cmac_dat459;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat460 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat460 <= ls2cmac_dat460;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat461 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat461 <= ls2cmac_dat461;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat462 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat462 <= ls2cmac_dat462;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat463 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat463 <= ls2cmac_dat463;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat464 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat464 <= ls2cmac_dat464;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat465 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat465 <= ls2cmac_dat465;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat466 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat466 <= ls2cmac_dat466;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat467 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat467 <= ls2cmac_dat467;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat468 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat468 <= ls2cmac_dat468;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat469 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat469 <= ls2cmac_dat469;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat470 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat470 <= ls2cmac_dat470;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat471 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat471 <= ls2cmac_dat471;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat472 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat472 <= ls2cmac_dat472;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat473 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat473 <= ls2cmac_dat473;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat474 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat474 <= ls2cmac_dat474;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat475 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat475 <= ls2cmac_dat475;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat476 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat476 <= ls2cmac_dat476;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat477 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat477 <= ls2cmac_dat477;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat478 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat478 <= ls2cmac_dat478;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat479 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat479 <= ls2cmac_dat479;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat480 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat480 <= ls2cmac_dat480;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat481 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat481 <= ls2cmac_dat481;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat482 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat482 <= ls2cmac_dat482;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat483 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat483 <= ls2cmac_dat483;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat484 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat484 <= ls2cmac_dat484;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat485 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat485 <= ls2cmac_dat485;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat486 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat486 <= ls2cmac_dat486;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat487 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat487 <= ls2cmac_dat487;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat488 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat488 <= ls2cmac_dat488;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat489 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat489 <= ls2cmac_dat489;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat490 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat490 <= ls2cmac_dat490;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat491 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat491 <= ls2cmac_dat491;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat492 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat492 <= ls2cmac_dat492;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat493 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat493 <= ls2cmac_dat493;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat494 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat494 <= ls2cmac_dat494;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat495 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat495 <= ls2cmac_dat495;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat496 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat496 <= ls2cmac_dat496;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat497 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat497 <= ls2cmac_dat497;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat498 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat498 <= ls2cmac_dat498;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat499 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat499 <= ls2cmac_dat499;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat500 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat500 <= ls2cmac_dat500;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat501 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat501 <= ls2cmac_dat501;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat502 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat502 <= ls2cmac_dat502;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat503 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat503 <= ls2cmac_dat503;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat504 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat504 <= ls2cmac_dat504;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat505 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat505 <= ls2cmac_dat505;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat506 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat506 <= ls2cmac_dat506;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat507 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat507 <= ls2cmac_dat507;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat508 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat508 <= ls2cmac_dat508;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat509 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat509 <= ls2cmac_dat509;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat510 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat510 <= ls2cmac_dat510;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat511 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat511 <= ls2cmac_dat511;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat512 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat512 <= ls2cmac_dat512;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat513 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat513 <= ls2cmac_dat513;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat514 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat514 <= ls2cmac_dat514;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat515 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat515 <= ls2cmac_dat515;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat516 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat516 <= ls2cmac_dat516;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat517 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat517 <= ls2cmac_dat517;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat518 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat518 <= ls2cmac_dat518;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat519 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat519 <= ls2cmac_dat519;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat520 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat520 <= ls2cmac_dat520;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat521 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat521 <= ls2cmac_dat521;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat522 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat522 <= ls2cmac_dat522;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat523 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat523 <= ls2cmac_dat523;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat524 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat524 <= ls2cmac_dat524;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat525 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat525 <= ls2cmac_dat525;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat526 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat526 <= ls2cmac_dat526;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat527 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat527 <= ls2cmac_dat527;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat528 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat528 <= ls2cmac_dat528;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat529 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat529 <= ls2cmac_dat529;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat530 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat530 <= ls2cmac_dat530;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat531 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat531 <= ls2cmac_dat531;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat532 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat532 <= ls2cmac_dat532;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat533 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat533 <= ls2cmac_dat533;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat534 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat534 <= ls2cmac_dat534;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat535 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat535 <= ls2cmac_dat535;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat536 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat536 <= ls2cmac_dat536;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat537 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat537 <= ls2cmac_dat537;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat538 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat538 <= ls2cmac_dat538;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat539 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat539 <= ls2cmac_dat539;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat540 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat540 <= ls2cmac_dat540;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat541 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat541 <= ls2cmac_dat541;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat542 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat542 <= ls2cmac_dat542;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat543 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat543 <= ls2cmac_dat543;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat544 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat544 <= ls2cmac_dat544;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat545 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat545 <= ls2cmac_dat545;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat546 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat546 <= ls2cmac_dat546;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat547 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat547 <= ls2cmac_dat547;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat548 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat548 <= ls2cmac_dat548;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat549 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat549 <= ls2cmac_dat549;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat550 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat550 <= ls2cmac_dat550;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat551 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat551 <= ls2cmac_dat551;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat552 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat552 <= ls2cmac_dat552;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat553 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat553 <= ls2cmac_dat553;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat554 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat554 <= ls2cmac_dat554;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat555 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat555 <= ls2cmac_dat555;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat556 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat556 <= ls2cmac_dat556;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat557 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat557 <= ls2cmac_dat557;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat558 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat558 <= ls2cmac_dat558;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat559 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat559 <= ls2cmac_dat559;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat560 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat560 <= ls2cmac_dat560;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat561 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat561 <= ls2cmac_dat561;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat562 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat562 <= ls2cmac_dat562;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat563 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat563 <= ls2cmac_dat563;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat564 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat564 <= ls2cmac_dat564;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat565 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat565 <= ls2cmac_dat565;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat566 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat566 <= ls2cmac_dat566;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat567 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat567 <= ls2cmac_dat567;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat568 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat568 <= ls2cmac_dat568;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat569 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat569 <= ls2cmac_dat569;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat570 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat570 <= ls2cmac_dat570;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat571 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat571 <= ls2cmac_dat571;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat572 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat572 <= ls2cmac_dat572;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat573 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat573 <= ls2cmac_dat573;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat574 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat574 <= ls2cmac_dat574;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat575 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat575 <= ls2cmac_dat575;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat576 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat576 <= ls2cmac_dat576;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat577 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat577 <= ls2cmac_dat577;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat578 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat578 <= ls2cmac_dat578;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat579 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat579 <= ls2cmac_dat579;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat580 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat580 <= ls2cmac_dat580;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat581 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat581 <= ls2cmac_dat581;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat582 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat582 <= ls2cmac_dat582;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat583 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat583 <= ls2cmac_dat583;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat584 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat584 <= ls2cmac_dat584;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat585 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat585 <= ls2cmac_dat585;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat586 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat586 <= ls2cmac_dat586;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat587 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat587 <= ls2cmac_dat587;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat588 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat588 <= ls2cmac_dat588;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat589 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat589 <= ls2cmac_dat589;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat590 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat590 <= ls2cmac_dat590;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat591 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat591 <= ls2cmac_dat591;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat592 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat592 <= ls2cmac_dat592;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat593 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat593 <= ls2cmac_dat593;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat594 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat594 <= ls2cmac_dat594;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat595 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat595 <= ls2cmac_dat595;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat596 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat596 <= ls2cmac_dat596;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat597 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat597 <= ls2cmac_dat597;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat598 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat598 <= ls2cmac_dat598;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat599 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat599 <= ls2cmac_dat599;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat600 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat600 <= ls2cmac_dat600;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat601 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat601 <= ls2cmac_dat601;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat602 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat602 <= ls2cmac_dat602;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat603 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat603 <= ls2cmac_dat603;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat604 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat604 <= ls2cmac_dat604;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat605 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat605 <= ls2cmac_dat605;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat606 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat606 <= ls2cmac_dat606;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat607 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat607 <= ls2cmac_dat607;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat608 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat608 <= ls2cmac_dat608;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat609 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat609 <= ls2cmac_dat609;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat610 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat610 <= ls2cmac_dat610;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat611 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat611 <= ls2cmac_dat611;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat612 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat612 <= ls2cmac_dat612;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat613 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat613 <= ls2cmac_dat613;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat614 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat614 <= ls2cmac_dat614;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat615 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat615 <= ls2cmac_dat615;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat616 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat616 <= ls2cmac_dat616;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat617 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat617 <= ls2cmac_dat617;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat618 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat618 <= ls2cmac_dat618;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat619 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat619 <= ls2cmac_dat619;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat620 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat620 <= ls2cmac_dat620;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat621 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat621 <= ls2cmac_dat621;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat622 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat622 <= ls2cmac_dat622;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat623 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat623 <= ls2cmac_dat623;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat624 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat624 <= ls2cmac_dat624;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat625 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat625 <= ls2cmac_dat625;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat626 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat626 <= ls2cmac_dat626;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat627 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat627 <= ls2cmac_dat627;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat628 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat628 <= ls2cmac_dat628;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat629 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat629 <= ls2cmac_dat629;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat630 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat630 <= ls2cmac_dat630;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat631 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat631 <= ls2cmac_dat631;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat632 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat632 <= ls2cmac_dat632;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat633 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat633 <= ls2cmac_dat633;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat634 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat634 <= ls2cmac_dat634;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat635 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat635 <= ls2cmac_dat635;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat636 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat636 <= ls2cmac_dat636;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat637 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat637 <= ls2cmac_dat637;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat638 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat638 <= ls2cmac_dat638;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat639 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat639 <= ls2cmac_dat639;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat640 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat640 <= ls2cmac_dat640;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat641 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat641 <= ls2cmac_dat641;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat642 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat642 <= ls2cmac_dat642;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat643 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat643 <= ls2cmac_dat643;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat644 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat644 <= ls2cmac_dat644;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat645 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat645 <= ls2cmac_dat645;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat646 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat646 <= ls2cmac_dat646;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat647 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat647 <= ls2cmac_dat647;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat648 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat648 <= ls2cmac_dat648;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat649 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat649 <= ls2cmac_dat649;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat650 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat650 <= ls2cmac_dat650;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat651 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat651 <= ls2cmac_dat651;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat652 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat652 <= ls2cmac_dat652;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat653 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat653 <= ls2cmac_dat653;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat654 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat654 <= ls2cmac_dat654;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat655 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat655 <= ls2cmac_dat655;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat656 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat656 <= ls2cmac_dat656;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat657 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat657 <= ls2cmac_dat657;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat658 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat658 <= ls2cmac_dat658;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat659 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat659 <= ls2cmac_dat659;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat660 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat660 <= ls2cmac_dat660;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat661 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat661 <= ls2cmac_dat661;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat662 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat662 <= ls2cmac_dat662;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat663 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat663 <= ls2cmac_dat663;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat664 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat664 <= ls2cmac_dat664;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat665 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat665 <= ls2cmac_dat665;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat666 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat666 <= ls2cmac_dat666;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat667 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat667 <= ls2cmac_dat667;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat668 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat668 <= ls2cmac_dat668;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat669 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat669 <= ls2cmac_dat669;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat670 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat670 <= ls2cmac_dat670;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat671 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat671 <= ls2cmac_dat671;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat672 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat672 <= ls2cmac_dat672;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat673 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat673 <= ls2cmac_dat673;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat674 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat674 <= ls2cmac_dat674;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat675 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat675 <= ls2cmac_dat675;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat676 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat676 <= ls2cmac_dat676;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat677 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat677 <= ls2cmac_dat677;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat678 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat678 <= ls2cmac_dat678;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat679 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat679 <= ls2cmac_dat679;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat680 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat680 <= ls2cmac_dat680;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat681 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat681 <= ls2cmac_dat681;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat682 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat682 <= ls2cmac_dat682;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat683 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat683 <= ls2cmac_dat683;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat684 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat684 <= ls2cmac_dat684;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat685 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat685 <= ls2cmac_dat685;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat686 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat686 <= ls2cmac_dat686;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat687 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat687 <= ls2cmac_dat687;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat688 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat688 <= ls2cmac_dat688;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat689 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat689 <= ls2cmac_dat689;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat690 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat690 <= ls2cmac_dat690;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat691 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat691 <= ls2cmac_dat691;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat692 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat692 <= ls2cmac_dat692;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat693 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat693 <= ls2cmac_dat693;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat694 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat694 <= ls2cmac_dat694;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat695 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat695 <= ls2cmac_dat695;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat696 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat696 <= ls2cmac_dat696;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat697 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat697 <= ls2cmac_dat697;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat698 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat698 <= ls2cmac_dat698;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat699 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat699 <= ls2cmac_dat699;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat700 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat700 <= ls2cmac_dat700;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat701 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat701 <= ls2cmac_dat701;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat702 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat702 <= ls2cmac_dat702;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat703 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat703 <= ls2cmac_dat703;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat704 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat704 <= ls2cmac_dat704;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat705 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat705 <= ls2cmac_dat705;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat706 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat706 <= ls2cmac_dat706;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat707 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat707 <= ls2cmac_dat707;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat708 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat708 <= ls2cmac_dat708;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat709 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat709 <= ls2cmac_dat709;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat710 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat710 <= ls2cmac_dat710;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat711 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat711 <= ls2cmac_dat711;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat712 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat712 <= ls2cmac_dat712;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat713 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat713 <= ls2cmac_dat713;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat714 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat714 <= ls2cmac_dat714;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat715 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat715 <= ls2cmac_dat715;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat716 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat716 <= ls2cmac_dat716;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat717 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat717 <= ls2cmac_dat717;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat718 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat718 <= ls2cmac_dat718;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat719 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat719 <= ls2cmac_dat719;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat720 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat720 <= ls2cmac_dat720;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat721 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat721 <= ls2cmac_dat721;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat722 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat722 <= ls2cmac_dat722;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat723 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat723 <= ls2cmac_dat723;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat724 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat724 <= ls2cmac_dat724;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat725 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat725 <= ls2cmac_dat725;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat726 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat726 <= ls2cmac_dat726;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat727 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat727 <= ls2cmac_dat727;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat728 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat728 <= ls2cmac_dat728;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat729 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat729 <= ls2cmac_dat729;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat730 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat730 <= ls2cmac_dat730;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat731 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat731 <= ls2cmac_dat731;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat732 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat732 <= ls2cmac_dat732;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat733 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat733 <= ls2cmac_dat733;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat734 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat734 <= ls2cmac_dat734;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat735 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat735 <= ls2cmac_dat735;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat736 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat736 <= ls2cmac_dat736;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat737 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat737 <= ls2cmac_dat737;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat738 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat738 <= ls2cmac_dat738;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat739 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat739 <= ls2cmac_dat739;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat740 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat740 <= ls2cmac_dat740;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat741 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat741 <= ls2cmac_dat741;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat742 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat742 <= ls2cmac_dat742;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat743 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat743 <= ls2cmac_dat743;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat744 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat744 <= ls2cmac_dat744;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat745 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat745 <= ls2cmac_dat745;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat746 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat746 <= ls2cmac_dat746;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat747 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat747 <= ls2cmac_dat747;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat748 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat748 <= ls2cmac_dat748;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat749 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat749 <= ls2cmac_dat749;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat750 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat750 <= ls2cmac_dat750;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat751 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat751 <= ls2cmac_dat751;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat752 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat752 <= ls2cmac_dat752;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat753 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat753 <= ls2cmac_dat753;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat754 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat754 <= ls2cmac_dat754;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat755 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat755 <= ls2cmac_dat755;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat756 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat756 <= ls2cmac_dat756;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat757 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat757 <= ls2cmac_dat757;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat758 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat758 <= ls2cmac_dat758;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat759 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat759 <= ls2cmac_dat759;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat760 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat760 <= ls2cmac_dat760;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat761 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat761 <= ls2cmac_dat761;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat762 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat762 <= ls2cmac_dat762;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat763 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat763 <= ls2cmac_dat763;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat764 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat764 <= ls2cmac_dat764;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat765 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat765 <= ls2cmac_dat765;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat766 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat766 <= ls2cmac_dat766;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat767 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat767 <= ls2cmac_dat767;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat768 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat768 <= ls2cmac_dat768;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat769 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat769 <= ls2cmac_dat769;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat770 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat770 <= ls2cmac_dat770;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat771 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat771 <= ls2cmac_dat771;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat772 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat772 <= ls2cmac_dat772;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat773 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat773 <= ls2cmac_dat773;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat774 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat774 <= ls2cmac_dat774;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat775 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat775 <= ls2cmac_dat775;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat776 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat776 <= ls2cmac_dat776;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat777 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat777 <= ls2cmac_dat777;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat778 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat778 <= ls2cmac_dat778;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat779 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat779 <= ls2cmac_dat779;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat780 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat780 <= ls2cmac_dat780;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat781 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat781 <= ls2cmac_dat781;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat782 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat782 <= ls2cmac_dat782;
        end
    end
    always_ff   @(posedge ytydla_conv_clk or negedge ytydla_core_rst_n) begin
        if (~ytydla_core_rst_n)begin
            conv_dat783 <= YTYDLA_DATA_LENGTH'b0;
        end
        else begin
            conv_dat783 <= ls2cmac_dat783;
        end
    end

    ytydla_conv_cmac cmac_0(
        .ytydla_core_clk    ytydla_core_clk,
        .ytydla_core_rst_n  ytydla_core_rst_n,
        .ls2cmac_dat0       ls2cmac_dat0,
        .ls2cmac_dat1       ls2cmac_dat1,
        .ls2cmac_dat2       ls2cmac_dat2,
        .ls2cmac_dat3       ls2cmac_dat3,
        .ls2cmac_dat4       ls2cmac_dat4,
        .ls2cmac_dat5       ls2cmac_dat5,
        .ls2cmac_dat6       ls2cmac_dat6,
        .ls2cmac_dat7       ls2cmac_dat7,
        .ls2cmac_dat8       ls2cmac_dat8,
        .ls2cmac_dat9       ls2cmac_dat9,
        .ls2cmac_dat10       ls2cmac_dat10,
        .ls2cmac_dat11       ls2cmac_dat11,
        .ls2cmac_dat12       ls2cmac_dat12,
        .ls2cmac_dat13       ls2cmac_dat13,
        .ls2cmac_dat14       ls2cmac_dat14,
        .ls2cmac_dat15       ls2cmac_dat15,
        .ls2cmac_dat16       ls2cmac_dat16,
        .ls2cmac_dat17       ls2cmac_dat17,
        .ls2cmac_dat18       ls2cmac_dat18,
        .ls2cmac_dat19       ls2cmac_dat19,
        .ls2cmac_dat20       ls2cmac_dat20,
        .ls2cmac_dat21       ls2cmac_dat21,
        .ls2cmac_dat22       ls2cmac_dat22,
        .ls2cmac_dat23       ls2cmac_dat23,
        .ls2cmac_dat24       ls2cmac_dat24,
        .ls2cmac_dat_bitmap  conv2cmac_dat_bitmap,
        .ls2cmac_wt0       ls2cmac_wt0,
        .ls2cmac_wt1       ls2cmac_wt1,
        .ls2cmac_wt2       ls2cmac_wt2,
        .ls2cmac_wt3       ls2cmac_wt3,
        .ls2cmac_wt4       ls2cmac_wt4,
        .ls2cmac_wt5       ls2cmac_wt5,
        .ls2cmac_wt6       ls2cmac_wt6,
        .ls2cmac_wt7       ls2cmac_wt7,
        .ls2cmac_wt8       ls2cmac_wt8,
        .ls2cmac_wt9       ls2cmac_wt9,
        .ls2cmac_wt10       ls2cmac_wt10,
        .ls2cmac_wt11       ls2cmac_wt11,
        .ls2cmac_wt12       ls2cmac_wt12,
        .ls2cmac_wt13       ls2cmac_wt13,
        .ls2cmac_wt14       ls2cmac_wt14,
        .ls2cmac_wt15       ls2cmac_wt15,
        .ls2cmac_wt16       ls2cmac_wt16,
        .ls2cmac_wt17       ls2cmac_wt17,
        .ls2cmac_wt18       ls2cmac_wt18,
        .ls2cmac_wt19       ls2cmac_wt19,
        .ls2cmac_wt20       ls2cmac_wt20,
        .ls2cmac_wt21       ls2cmac_wt21,
        .ls2cmac_wt22       ls2cmac_wt22,
        .ls2cmac_wt23       ls2cmac_wt23,
        .ls2cmac_wt24       ls2cmac_wt24,
        .ls2cmac_wt_bitmap  conv2cmac_wt_bitmap);
    

endmodule
