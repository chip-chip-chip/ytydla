// ytydla_define.svh


`define YTYDLA_DATA_LENGTH  32
`define YTYDLA_DATA_DOTPOT  12
